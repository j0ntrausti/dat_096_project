


-- This is a Linear phase FIR filter of type 1. Has N coeff. and N-1 inputs.
-- The filter is written GENERIC so it is defined as;
--                            WIDTH = number of bits
--                            N = number of tabs   
--			      M = Channel filter type, (to maximise the available space for multiplication)
-- Takes in, GENERIC values WIDTH (nr. of bits), N number of tabs, x[n].
-- Sends out finihs signal, and y[n] (note double size, need to take the 12 last bits)
-- Authors: Jo³n Trausti
library ieee;
use ieee.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

entity Block_Filter_250 is
    GENERIC(WIDTH    :integer     :=12;
        N :integer    :=188);
    PORT(    reset:IN STD_LOGIC;
           clk:IN STD_LOGIC;
           clk312K:IN STD_LOGIC;
           clk625K:IN STD_LOGIC;
           x:IN signed(WIDTH-1 DOWNTO 0);
           y:OUT signed(WIDTH-1 DOWNTO 0);
           finished:OUT STD_LOGIC);
end Block_Filter_250;



architecture behaiv_arch of Block_Filter_250 is


-- New signals
signal i    :integer range 0 to N+3; --index for how many clkcykles the calculation have been running
signal finished_sig,GoOn,Load_On    :STD_LOGIC :='0';
signal a_s,b_s    :signed(2*WIDTH-1 downto 0);--temporary output
signal x_sig :signed(WIDTH-1 downto 0);

type a_pipe is array (0 to N-1) of signed(WIDTH-1 downto 0);
type a_queue2multi is array (0 to N-1) of signed(WIDTH-1 downto 0);
type a_tL is array (0 to N-1) of signed(WIDTH-1 downto 0);

signal pipe    		: a_pipe;
signal queue2multi	:a_queue2multi;
signal t		:a_tL;




-- Old signals



begin


--x_sig(WIDTH-1 downto 4) <= x;
--x_sig(3 downto 0) <= (others => '0');
process(clk,reset)
begin

    -- This will set all the x's to zero, resetting everything.
    -- so when the program start all values have zeros except for the coefficients
    if(reset='1') then
        i<=0;    -- reset the counter
        a_s <= (others => '0');
	b_s <= (others => '0');
        y <= (others => '0');
        finished <= '0';
        finished_sig <= '1';
        for i in 0 to (N-1) loop
               pipe(i)<=(others=> '0');
               queue2multi(i)<=(others=> '0');
        end loop;
        

        -- here the coeff. comes in for ex.
t(0)<="0000000000111011";
        t(1)<="0000000010100010";
        t(2)<="0000000011111111";
        t(3)<="0000000011110100";
        t(4)<="0000000001011011";
        t(5)<="1111111110001000";
        t(6)<="1111111100010000";
        t(7)<="1111111101000001";
        t(8)<="1111111111010000";
        t(9)<="0000000000100011";
        t(10)<="1111111111110000";
        t(11)<="1111111110000111";
        t(12)<="1111111101101101";
        t(13)<="1111111110111101";
        t(14)<="0000000000010010";
        t(15)<="0000000000000101";
        t(16)<="1111111110110001";
        t(17)<="1111111110001001";
        t(18)<="1111111111000011";
        t(19)<="0000000000010101";
        t(20)<="0000000000010100";
        t(21)<="1111111111000110";
        t(22)<="1111111110010110";
        t(23)<="1111111111001001";
        t(24)<="0000000000011101";
        t(25)<="0000000000100011";
        t(26)<="1111111111010011";
        t(27)<="1111111110011011";
        t(28)<="1111111111001011";
        t(29)<="0000000000100111";
        t(30)<="0000000000110010";
        t(31)<="1111111111011100";
        t(32)<="1111111110011010";
        t(33)<="1111111111001010";
        t(34)<="0000000000110000";
        t(35)<="0000000001000010";
        t(36)<="1111111111100101";
        t(37)<="1111111110010101";
        t(38)<="1111111111000100";
        t(39)<="0000000000111000";
        t(40)<="0000000001010100";
        t(41)<="1111111111101101";
        t(42)<="1111111110001100";
        t(43)<="1111111110111011";
        t(44)<="0000000001000000";
        t(45)<="0000000001100111";
        t(46)<="1111111111110101";
        t(47)<="1111111110000001";
        t(48)<="1111111110101110";
        t(49)<="0000000001000110";
        t(50)<="0000000001111100";
        t(51)<="1111111111111111";
        t(52)<="1111111101110100";
        t(53)<="1111111110011101";
        t(54)<="0000000001001100";
        t(55)<="0000000010010100";
        t(56)<="0000000000001010";
        t(57)<="1111111101100100";
        t(58)<="1111111110001000";
        t(59)<="0000000001010001";
        t(60)<="0000000010110000";
        t(61)<="0000000000011000";
        t(62)<="1111111101010000";
        t(63)<="1111111101101110";
        t(64)<="0000000001010110";
        t(65)<="0000000011010001";
        t(66)<="0000000000101010";
        t(67)<="1111111100111001";
        t(68)<="1111111101001101";
        t(69)<="0000000001011010";
        t(70)<="0000000011111001";
        t(71)<="0000000001000001";
        t(72)<="1111111100011101";
        t(73)<="1111111100100010";
        t(74)<="0000000001011110";
        t(75)<="0000000100101011";
        t(76)<="0000000001011110";
        t(77)<="1111111011111001";
        t(78)<="1111111011101001";
        t(79)<="0000000001100001";
        t(80)<="0000000101101110";
        t(81)<="0000000010001000";
        t(82)<="1111111011001001";
        t(83)<="1111111010011001";
        t(84)<="0000000001100100";
        t(85)<="0000000111001101";
        t(86)<="0000000011000110";
        t(87)<="1111111010000011";
        t(88)<="1111111000100001";
        t(89)<="0000000001100110";
        t(90)<="0000001001100000";
        t(91)<="0000000100101001";
        t(92)<="1111111000010001";
        t(93)<="1111110101010100";
        t(94)<="0000000001101000";
        t(95)<="0000001101101101";
        t(96)<="0000000111101000";
        t(97)<="1111110100101101";
        t(98)<="1111101110011101";
        t(99)<="0000000001101001";
        t(100)<="0000011000001100";
        t(101)<="0000001111111111";
        t(102)<="1111101001011011";
        t(103)<="1111010100010011";
        t(104)<="0000000001101001";
        t(105)<="0001100111110011";
        t(106)<="0010111110001110";
        t(107)<="0010111110001110";
        t(108)<="0001100111110011";
        t(109)<="0000000001101001";
        t(110)<="1111010100010011";
        t(111)<="1111101001011011";
        t(112)<="0000001111111111";
        t(113)<="0000011000001100";
        t(114)<="0000000001101001";
        t(115)<="1111101110011101";
        t(116)<="1111110100101101";
        t(117)<="0000000111101000";
        t(118)<="0000001101101101";
        t(119)<="0000000001101000";
        t(120)<="1111110101010100";
        t(121)<="1111111000010001";
        t(122)<="0000000100101001";
        t(123)<="0000001001100000";
        t(124)<="0000000001100110";
        t(125)<="1111111000100001";
        t(126)<="1111111010000011";
        t(127)<="0000000011000110";
        t(128)<="0000000111001101";
        t(129)<="0000000001100100";
        t(130)<="1111111010011001";
        t(131)<="1111111011001001";
        t(132)<="0000000010001000";
        t(133)<="0000000101101110";
        t(134)<="0000000001100001";
        t(135)<="1111111011101001";
        t(136)<="1111111011111001";
        t(137)<="0000000001011110";
        t(138)<="0000000100101011";
        t(139)<="0000000001011110";
        t(140)<="1111111100100010";
        t(141)<="1111111100011101";
        t(142)<="0000000001000001";
        t(143)<="0000000011111001";
        t(144)<="0000000001011010";
        t(145)<="1111111101001101";
        t(146)<="1111111100111001";
        t(147)<="0000000000101010";
        t(148)<="0000000011010001";
        t(149)<="0000000001010110";
        t(150)<="1111111101101110";
        t(151)<="1111111101010000";
        t(152)<="0000000000011000";
        t(153)<="0000000010110000";
        t(154)<="0000000001010001";
        t(155)<="1111111110001000";
        t(156)<="1111111101100100";
        t(157)<="0000000000001010";
        t(158)<="0000000010010100";
        t(159)<="0000000001001100";
        t(160)<="1111111110011101";
        t(161)<="1111111101110100";
        t(162)<="1111111111111111";
        t(163)<="0000000001111100";
        t(164)<="0000000001000110";
        t(165)<="1111111110101110";
        t(166)<="1111111110000001";
        t(167)<="1111111111110101";
        t(168)<="0000000001100111";
        t(169)<="0000000001000000";
        t(170)<="1111111110111011";
        t(171)<="1111111110001100";
        t(172)<="1111111111101101";
        t(173)<="0000000001010100";
        t(174)<="0000000000111000";
        t(175)<="1111111111000100";
        t(176)<="1111111110010101";
        t(177)<="1111111111100101";
        t(178)<="0000000001000010";
        t(179)<="0000000000110000";
        t(180)<="1111111111001010";
        t(181)<="1111111110011010";
        t(182)<="1111111111011100";
        t(183)<="0000000000110010";
        t(184)<="0000000000100111";
        t(185)<="1111111111001011";
        t(186)<="1111111110011011";
        t(187)<="1111111111010011";
        t(188)<="0000000000100011";
        t(189)<="0000000000011101";
        t(190)<="1111111111001001";
        t(191)<="1111111110010110";
        t(192)<="1111111111000110";
        t(193)<="0000000000010100";
        t(194)<="0000000000010101";
        t(195)<="1111111111000011";
        t(196)<="1111111110001001";
        t(197)<="1111111110110001";
        t(198)<="0000000000000101";
        t(199)<="0000000000010010";
        t(200)<="1111111110111101";
        t(201)<="1111111101101101";
        t(202)<="1111111110000111";
        t(203)<="1111111111110000";
        t(204)<="0000000000100011";
        t(205)<="1111111111010000";
        t(206)<="1111111101000001";
        t(207)<="1111111100010000";
        t(208)<="1111111110001000";
        t(209)<="0000000001011011";
        t(210)<="0000000011110100";
        t(211)<="0000000011111111";
        t(212)<="0000000010100010";
        t(213)<="0000000000111011";






    elsif (rising_edge(clk)) then
--------------------------------------------------------------------    
-----------------------------SENDING OUT ---------------------------    
--------------------------------------------------------------------       
        if(clk312K = '1') then   
		Load_On<='1';
        	a_s <= (others => '0');
        	b_s <= (others => '0');
            	finished_sig <= '0';
           	finished<='0';
         	i<=0;
	elsif(finished_sig = '0' AND Load_On='0' AND GoOn='1') then
		if(i<N/2) then
			a_s <= a_s + (queue2multi(2*i)*t(2*i));
			b_s <= b_s + (queue2multi(2*i+1)*t(2*i+1));
			i <= i+1;
		else
			finished <= '1';
                	finished_sig <= '1';
               		y <= a_s(2*WIDTH-2 downto WIDTH-1) + b_s(2*WIDTH-2 downto WIDTH-1);
		end if;
		
        end if;
--------------------------------------------------------------------    
-----------------------------READING IN ----------------------------    
--------------------------------------------------------------------  

	if (clk625K='1' ) then 
		pipe <= signed(x)&pipe(0 to pipe'length-2);
	elsif(Load_On ='1') then
		for j in 0 to N-1 loop
             	   queue2multi(j)<= pipe(j);
         	end loop;
		GoOn<='1';  
		Load_On<='0';
	end if;

    end if;
end process;

end behaiv_arch;
