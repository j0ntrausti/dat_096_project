

-- This is a Linear phase FIR filter of type 1. Has N coeff. and N-1 inputs.
-- The filter is written generic so it is defined as;
--                            Width = number of bits
--                            N = number of tabs   
--			      M = Channel filter type, (to maximise the available space for multiplication)
-- Takes in, generic values width (nr. of bits), N number of tabs, x[n].
-- Sends out finihs signal, and y[n] (note double size, need to take the 12 last bits)
-- Authors: Jo³n Trausti
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity FastFilter is
    generic(Width    :integer     :=24;
        N :integer    :=20);
	--M :integer :=0);
    port(    reset:IN STD_LOGIC;
           clk:IN STD_LOGIC;
           clk250k:IN STD_LOGIC;
           clk6M:IN STD_LOGIC;
           x:IN signed(width-13 DOWNTO 0);
           y:OUT signed(WIDTH-13 DOWNTO 0);
           finished:OUT STD_LOGIC);
end FastFilter;



architecture behaiv_arch of FastFilter is


-- New signals
signal swapping    :std_logic :='0'; --this shall trigger when start goes to '1' and go down when start goes to '0' to see if there is a new x or not
signal i    :integer range 0 to N+3; --index for how many clkcykles the calculation have been running

signal finished_sig,GoOn,Load_On   :std_logic :='0';
signal a_s,b_s,c_s,d_s,e_s,f_s     :signed(2*width-1 downto 0);--temporary output
signal x_sig                       :signed(width-1 downto 0);


type a_array is array (0 to (N-1)) of signed(width-1 downto 0);

signal t		:a_array;
signal queue2multi	:a_array;
signal pipe		:a_array;



-- Old signals



begin

x_sig(width-1 downto 12) <= x;
x_sig(11 downto 0) <= (others => '0');

process(clk,reset)
begin

    -- This will set all the x's to zero, resetting everything.
    -- so when the program start all values have zeros except for the coefficients
    if(reset='1') then
        i<=0;    -- reset the counte
        y <= (others => '0');
        finished <= '0';
        finished_sig <= '1';
	a_s <= (others => '0');
        b_s <= (others => '0');
        c_s <= (others => '0');
        d_s <= (others => '0');
        e_s <= (others => '0');
	f_s <= (others => '0');
        for i in 0 to (N-1) loop
               pipe(i)<=(others=> '0');
               queue2multi(i)<=(others=> '0');
        end loop;
        

        -- here the coeff. comes in for ex.

		



t(0)<="111111111111111111111111";
t(1)<="111111111111010010101011";
t(2)<="111111111111101111000100";
t(3)<="111111111111101010011100";
t(4)<="111111111111100110110001";
t(5)<="111111111111100010110000";
t(6)<="111111111111011110011110";
t(7)<="111111111111011001111001";
t(8)<="111111111111010101000101";
t(9)<="111111111111010000000010";
t(10)<="111111111111001010110010";
t(11)<="111111111111000101010110";
t(12)<="111111111110111111110001";
t(13)<="111111111110111010000101";
t(14)<="111111111110110100010101";
t(15)<="111111111110101110100100";
t(16)<="111111111110101000110100";
t(17)<="111111111110100011001001";
t(18)<="111111111110011101100110";
t(19)<="111111111110011000001101";
t(20)<="111111111110010011000011";
t(21)<="111111111110001110001001";
t(22)<="111111111110001001100101";
t(23)<="111111111110000101011001";
t(24)<="111111111110000001101001";
t(25)<="111111111101111110010110";
t(26)<="111111111101111011100110";
t(27)<="111111111101111001011001";
t(28)<="111111111101110111110011";
t(29)<="111111111101110110110100";
t(30)<="111111111101110110100000";
t(31)<="111111111101110110110110";
t(32)<="111111111101110111111011";
t(33)<="111111111101111001101100";
t(34)<="111111111101111100001100";
t(35)<="111111111101111111010111";
t(36)<="111111111110000011001111";
t(37)<="111111111110000111110010";
t(38)<="111111111110001101000010";
t(39)<="111111111110010010111000";
t(40)<="111111111110011001010100";
t(41)<="111111111110100000010001";
t(42)<="111111111110100111101111";
t(43)<="111111111110101111101001";
t(44)<="111111111110110111111011";
t(45)<="111111111111000000011101";
t(46)<="111111111111001001010100";
t(47)<="111111111111010010010011";
t(48)<="111111111111011011010101";
t(49)<="111111111111100100011011";
t(50)<="111111111111101101011010";
t(51)<="111111111111111111111111";
t(52)<="111111111111111111111111";
t(53)<="000000000000000111001110";
t(54)<="000000000000001111001010";
t(55)<="000000000000010110101010";
t(56)<="000000000000011101101010";
t(57)<="000000000000100100000100";
t(58)<="000000000000101001110111";
t(59)<="000000000000101110111111";
t(60)<="000000000000110011011001";
t(61)<="000000000000110111000011";
t(62)<="000000000000111001111100";
t(63)<="000000000000111100000010";
t(64)<="000000000000111101010110";
t(65)<="000000000000111101110111";
t(66)<="000000000000111101100101";
t(67)<="000000000000111100100011";
t(68)<="000000000000111010110010";
t(69)<="000000000000111000010011";
t(70)<="000000000000110101001011";
t(71)<="000000000000110001011011";
t(72)<="000000000000101101001001";
t(73)<="000000000000101000011000";
t(74)<="000000000000100011001100";
t(75)<="000000000000011101101010";
t(76)<="000000000000010111110111";
t(77)<="000000000000010001111000";
t(78)<="000000000000001011110010";
t(79)<="000000000000000101101011";
t(80)<="111111111111111111111111";
t(81)<="111111111111111111111111";
t(82)<="111111111111111111111111";
t(83)<="111111111111101110100011";
t(84)<="111111111111101001011111";
t(85)<="111111111111100100110100";
t(86)<="111111111111100000101000";
t(87)<="111111111111011100111101";
t(88)<="111111111111011001110111";
t(89)<="111111111111010111010110";
t(90)<="111111111111010101011110";
t(91)<="111111111111010100001110";
t(92)<="111111111111010011101000";
t(93)<="111111111111010011101100";
t(94)<="111111111111010100011001";
t(95)<="111111111111010101101101";
t(96)<="111111111111010111100111";
t(97)<="111111111111011010000101";
t(98)<="111111111111011101000100";
t(99)<="111111111111100000100001";
t(100)<="111111111111100100011000";
t(101)<="111111111111101000100101";
t(102)<="111111111111101101000101";
t(103)<="111111111111110001110011";
t(104)<="111111111111111111111111";
t(105)<="111111111111111111111111";
t(106)<="000000000000000000100000";
t(107)<="000000000000000101010110";
t(108)<="000000000000001010000100";
t(109)<="000000000000001110100011";
t(110)<="000000000000010010110001";
t(111)<="000000000000010110101001";
t(112)<="000000000000011010001001";
t(113)<="000000000000011101001011";
t(114)<="000000000000011111110000";
t(115)<="000000000000100001110011";
t(116)<="000000000000100011010100";
t(117)<="000000000000100100010001";
t(118)<="000000000000100100101010";
t(119)<="000000000000100100011110";
t(120)<="000000000000100011101111";
t(121)<="000000000000100010011100";
t(122)<="000000000000100000101000";
t(123)<="000000000000011110010101";
t(124)<="000000000000011011100110";
t(125)<="000000000000011000011100";
t(126)<="000000000000010100111100";
t(127)<="000000000000010001001000";
t(128)<="000000000000001101000110";
t(129)<="000000000000001000111001";
t(130)<="000000000000000100100110";
t(131)<="000000000000000000010000";
t(132)<="111111111111111111111111";
t(133)<="111111111111111111111111";
t(134)<="111111111111111111111111";
t(135)<="111111111111101111110110";
t(136)<="111111111111101100010011";
t(137)<="111111111111101001000110";
t(138)<="111111111111100110010001";
t(139)<="111111111111100011111000";
t(140)<="111111111111100001111101";
t(141)<="111111111111100000100000";
t(142)<="111111111111011111100101";
t(143)<="111111111111011111001011";
t(144)<="111111111111011111010011";
t(145)<="111111111111011111111011";
t(146)<="111111111111100001000101";
t(147)<="111111111111100010101110";
t(148)<="111111111111100100110100";
t(149)<="111111111111100111010110";
t(150)<="111111111111101010010000";
t(151)<="111111111111101101011111";
t(152)<="111111111111110001000001";
t(153)<="111111111111111111111111";
t(154)<="111111111111111111111111";
t(155)<="111111111111111111111111";
t(156)<="000000000000000000101111";
t(157)<="000000000000000100110000";
t(158)<="000000000000001000101100";
t(159)<="000000000000001100011101";
t(160)<="000000000000010000000001";
t(161)<="000000000000010011010011";
t(162)<="000000000000010110010001";
t(163)<="000000000000011000110111";
t(164)<="000000000000011011000010";
t(165)<="000000000000011100110001";
t(166)<="000000000000011110000010";
t(167)<="000000000000011110110011";
t(168)<="000000000000011111000100";
t(169)<="000000000000011110110101";
t(170)<="000000000000011110000101";
t(171)<="000000000000011100110111";
t(172)<="000000000000011011001010";
t(173)<="000000000000011001000001";
t(174)<="000000000000010110011111";
t(175)<="000000000000010011100101";
t(176)<="000000000000010000010111";
t(177)<="000000000000001100111000";
t(178)<="000000000000001001001101";
t(179)<="000000000000000101010111";
t(180)<="000000000000000001011101";
t(181)<="111111111111111111111111";
t(182)<="111111111111111111111111";
t(183)<="111111111111111111111111";
t(184)<="111111111111110010010000";
t(185)<="111111111111101110111000";
t(186)<="111111111111101011110010";
t(187)<="111111111111101001000001";
t(188)<="111111111111100110101001";
t(189)<="111111111111100100101011";
t(190)<="111111111111100011001010";
t(191)<="111111111111100010000111";
t(192)<="111111111111100001100100";
t(193)<="111111111111100001100001";
t(194)<="111111111111100001111110";
t(195)<="111111111111100010111011";
t(196)<="111111111111100100010110";
t(197)<="111111111111100110001111";
t(198)<="111111111111101000100010";
t(199)<="111111111111101011001111";
t(200)<="111111111111101110010001";
t(201)<="111111111111110001100110";
t(202)<="111111111111111111111111";
t(203)<="111111111111111111111111";
t(204)<="111111111111111111111111";
t(205)<="000000000000000000101110";
t(206)<="000000000000000100101001";
t(207)<="000000000000001000011111";
t(208)<="000000000000001100001101";
t(209)<="000000000000001111101101";
t(210)<="000000000000010010111110";
t(211)<="000000000000010101111010";
t(212)<="000000000000011000100000";
t(213)<="000000000000011010101100";
t(214)<="000000000000011100011100";
t(215)<="000000000000011101101101";
t(216)<="000000000000011110100000";
t(217)<="000000000000011110110010";
t(218)<="000000000000011110100100";
t(219)<="000000000000011101110101";
t(220)<="000000000000011100100111";
t(221)<="000000000000011010111010";
t(222)<="000000000000011000110001";
t(223)<="000000000000010110001100";
t(224)<="000000000000010011010001";
t(225)<="000000000000010000000000";
t(226)<="000000000000001100011110";
t(227)<="000000000000001000101110";
t(228)<="000000000000000100110100";
t(229)<="000000000000000000110101";
t(230)<="111111111111111111111111";
t(231)<="111111111111111111111111";
t(232)<="111111111111111111111111";
t(233)<="111111111111110001010010";
t(234)<="111111111111101101110101";
t(235)<="111111111111101010101011";
t(236)<="111111111111100111110111";
t(237)<="111111111111100101011011";
t(238)<="111111111111100011011100";
t(239)<="111111111111100001111011";
t(240)<="111111111111100000111001";
t(241)<="111111111111100000011000";
t(242)<="111111111111100000011001";
t(243)<="111111111111100000111011";
t(244)<="111111111111100001111110";
t(245)<="111111111111100011100010";
t(246)<="111111111111100101100100";
t(247)<="111111111111101000000010";
t(248)<="111111111111101010111011";
t(249)<="111111111111101110001010";
t(250)<="111111111111110001101101";
t(251)<="111111111111111111111111";
t(252)<="111111111111111111111111";
t(253)<="111111111111111111111111";
t(254)<="000000000000000001110001";
t(255)<="000000000000000101111010";
t(256)<="000000000000001001111110";
t(257)<="000000000000001101111000";
t(258)<="000000000000010001100101";
t(259)<="000000000000010100111111";
t(260)<="000000000000011000000100";
t(261)<="000000000000011010110001";
t(262)<="000000000000011101000001";
t(263)<="000000000000011110110011";
t(264)<="000000000000100000000101";
t(265)<="000000000000100000110101";
t(266)<="000000000000100001000010";
t(267)<="000000000000100000101100";
t(268)<="000000000000011111110100";
t(269)<="000000000000011110011001";
t(270)<="000000000000011100011110";
t(271)<="000000000000011010000011";
t(272)<="000000000000010111001101";
t(273)<="000000000000010011111101";
t(274)<="000000000000010000010111";
t(275)<="000000000000001100011111";
t(276)<="000000000000001000011000";
t(277)<="000000000000000100001000";
t(278)<="111111111111111111111111";
t(279)<="111111111111111111111111";
t(280)<="111111111111111111111111";
t(281)<="111111111111111111111111";
t(282)<="111111111111101110111110";
t(283)<="111111111111101011010001";
t(284)<="111111111111100111111001";
t(285)<="111111111111100100111010";
t(286)<="111111111111100010010111";
t(287)<="111111111111100000010010";
t(288)<="111111111111011110101111";
t(289)<="111111111111011101101111";
t(290)<="111111111111011101010011";
t(291)<="111111111111011101011011";
t(292)<="111111111111011110001001";
t(293)<="111111111111011111011011";
t(294)<="111111111111100001010000";
t(295)<="111111111111100011100110";
t(296)<="111111111111100110011011";
t(297)<="111111111111101001101100";
t(298)<="111111111111101101010110";
t(299)<="111111111111110001010101";
t(300)<="111111111111111111111111";
t(301)<="111111111111111111111111";
t(302)<="111111111111111111111111";
t(303)<="000000000000000011001011";
t(304)<="000000000000000111110000";
t(305)<="000000000000001100001110";
t(306)<="000000000000010000100000";
t(307)<="000000000000010100100010";
t(308)<="000000000000011000001111";
t(309)<="000000000000011011100100";
t(310)<="000000000000011110011100";
t(311)<="000000000000100000110101";
t(312)<="000000000000100010101011";
t(313)<="000000000000100011111101";
t(314)<="000000000000100100101010";
t(315)<="000000000000100100101111";
t(316)<="000000000000100100001101";
t(317)<="000000000000100011000101";
t(318)<="000000000000100001010111";
t(319)<="000000000000011111000101";
t(320)<="000000000000011100010001";
t(321)<="000000000000011000111110";
t(322)<="000000000000010101001111";
t(323)<="000000000000010001001000";
t(324)<="000000000000001100101111";
t(325)<="000000000000001000000101";
t(326)<="000000000000000011010010";
t(327)<="111111111111111111111111";
t(328)<="111111111111111111111111";
t(329)<="111111111111111111111111";
t(330)<="111111111111110000000111";
t(331)<="111111111111101011101110";
t(332)<="111111111111100111101001";
t(333)<="111111111111100011111101";
t(334)<="111111111111100000101101";
t(335)<="111111111111011101111110";
t(336)<="111111111111011011110010";
t(337)<="111111111111011010001100";
t(338)<="111111111111011001001101";
t(339)<="111111111111011000111000";
t(340)<="111111111111011001001100";
t(341)<="111111111111011010001001";
t(342)<="111111111111011011101111";
t(343)<="111111111111011101111100";
t(344)<="111111111111100000101111";
t(345)<="111111111111100100000011";
t(346)<="111111111111100111110110";
t(347)<="111111111111101100000101";
t(348)<="111111111111110000101001";
t(349)<="111111111111111111111111";
t(350)<="111111111111111111111111";
t(351)<="111111111111111111111111";
t(352)<="000000000000000100111100";
t(353)<="000000000000001010000101";
t(354)<="000000000000001111000110";
t(355)<="000000000000010011111000";
t(356)<="000000000000011000010111";
t(357)<="000000000000011100011101";
t(358)<="000000000000100000000110";
t(359)<="000000000000100011001111";
t(360)<="000000000000100101110011";
t(361)<="000000000000100111101111";
t(362)<="000000000000101001000010";
t(363)<="000000000000101001101001";
t(364)<="000000000000101001100101";
t(365)<="000000000000101000110100";
t(366)<="000000000000100111010111";
t(367)<="000000000000100101010000";
t(368)<="000000000000100010100000";
t(369)<="000000000000011111001011";
t(370)<="000000000000011011010011";
t(371)<="000000000000010110111101";
t(372)<="000000000000010010001101";
t(373)<="000000000000001101001000";
t(374)<="000000000000000111110011";
t(375)<="000000000000000010010100";
t(376)<="111111111111111111111111";
t(377)<="111111111111111111111111";
t(378)<="111111111111110001110100";
t(379)<="111111111111101100100110";
t(380)<="111111111111100111101100";
t(381)<="111111111111100011001001";
t(382)<="111111111111011111000100";
t(383)<="111111111111011011100000";
t(384)<="111111111111011000100010";
t(385)<="111111111111010110001101";
t(386)<="111111111111010100100100";
t(387)<="111111111111010011101001";
t(388)<="111111111111010011011100";
t(389)<="111111111111010011111111";
t(390)<="111111111111010101010001";
t(391)<="111111111111010111010001";
t(392)<="111111111111011001111101";
t(393)<="111111111111011101010010";
t(394)<="111111111111100001001110";
t(395)<="111111111111100101101100";
t(396)<="111111111111101010101000";
t(397)<="111111111111101111111100";
t(398)<="111111111111111111111111";
t(399)<="111111111111111111111111";
t(400)<="000000000000000001010100";
t(401)<="000000000000000111010000";
t(402)<="000000000000001101000111";
t(403)<="000000000000010010110001";
t(404)<="000000000000011000001011";
t(405)<="000000000000011101001100";
t(406)<="000000000000100001110000";
t(407)<="000000000000100101110001";
t(408)<="000000000000101001001100";
t(409)<="000000000000101011111100";
t(410)<="000000000000101101111111";
t(411)<="000000000000101111010001";
t(412)<="000000000000101111110001";
t(413)<="000000000000101111011110";
t(414)<="000000000000101110011001";
t(415)<="000000000000101100100010";
t(416)<="000000000000101001111011";
t(417)<="000000000000100110100110";
t(418)<="000000000000100010100111";
t(419)<="000000000000011110000001";
t(420)<="000000000000011000111010";
t(421)<="000000000000010011010110";
t(422)<="000000000000001101011100";
t(423)<="000000000000000111010001";
t(424)<="000000000000000000111100";
t(425)<="111111111111111111111111";
t(426)<="111111111111111111111111";
t(427)<="111111111111101110000100";
t(428)<="111111111111101000001010";
t(429)<="111111111111100010100111";
t(430)<="111111111111011101100001";
t(431)<="111111111111011000111111";
t(432)<="111111111111010101000100";
t(433)<="111111111111010001110101";
t(434)<="111111111111001111010111";
t(435)<="111111111111001101101011";
t(436)<="111111111111001100110100";
t(437)<="111111111111001100110100";
t(438)<="111111111111001101101010";
t(439)<="111111111111001111010110";
t(440)<="111111111111010001110111";
t(441)<="111111111111010101001001";
t(442)<="111111111111011001001011";
t(443)<="111111111111011101110111";
t(444)<="111111111111100011001010";
t(445)<="111111111111101000111101";
t(446)<="111111111111101111001011";
t(447)<="111111111111111111111111";
t(448)<="111111111111111111111111";
t(449)<="000000000000000011010100";
t(450)<="000000000000001010001001";
t(451)<="000000000000010000110110";
t(452)<="000000000000010111010011";
t(453)<="000000000000011101011010";
t(454)<="000000000000100011000100";
t(455)<="000000000000101000001011";
t(456)<="000000000000101100101001";
t(457)<="000000000000110000011001";
t(458)<="000000000000110011010111";
t(459)<="000000000000110101100000";
t(460)<="000000000000110110110000";
t(461)<="000000000000110111000110";
t(462)<="000000000000110110100001";
t(463)<="000000000000110101000011";
t(464)<="000000000000110010101011";
t(465)<="000000000000101111011100";
t(466)<="000000000000101011011001";
t(467)<="000000000000100110100111";
t(468)<="000000000000100001001001";
t(469)<="000000000000011011000111";
t(470)<="000000000000010100100100";
t(471)<="000000000000001101101010";
t(472)<="000000000000000110011110";
t(473)<="111111111111111111111111";
t(474)<="111111111111111111111111";
t(475)<="111111111111110000100000";
t(476)<="111111111111101001011100";
t(477)<="111111111111100010101101";
t(478)<="111111111111011100011100";
t(479)<="111111111111010110101101";
t(480)<="111111111111010001101001";
t(481)<="111111111111001101010011";
t(482)<="111111111111001001110010";
t(483)<="111111111111000111001010";
t(484)<="111111111111000101011101";
t(485)<="111111111111000100101110";
t(486)<="111111111111000100111110";
t(487)<="111111111111000110001100";
t(488)<="111111111111001000011001";
t(489)<="111111111111001011100010";
t(490)<="111111111111001111100100";
t(491)<="111111111111010100011011";
t(492)<="111111111111011010000011";
t(493)<="111111111111100000010101";
t(494)<="111111111111100111001011";
t(495)<="111111111111101110011111";
t(496)<="111111111111111111111111";
t(497)<="111111111111111111111111";
t(498)<="000000000000000101111010";
t(499)<="000000000000001101110010";
t(500)<="000000000000010101011111";
t(501)<="000000000000011100111000";
t(502)<="000000000000100011110101";
t(503)<="000000000000101010001110";
t(504)<="000000000000101111111101";
t(505)<="000000000000110100111011";
t(506)<="000000000000111001000010";
t(507)<="000000000000111100001111";
t(508)<="000000000000111110011100";
t(509)<="000000000000111111100111";
t(510)<="000000000000111111110000";
t(511)<="000000000000111110110100";
t(512)<="000000000000111100110101";
t(513)<="000000000000111001110100";
t(514)<="000000000000110101110100";
t(515)<="000000000000110000111001";
t(516)<="000000000000101011001001";
t(517)<="000000000000100100100111";
t(518)<="000000000000011101011101";
t(519)<="000000000000010101110000";
t(520)<="000000000000001101101000";
t(521)<="000000000000000101001111";
t(522)<="111111111111111111111111";
t(523)<="111111111111111111111111";
t(524)<="111111111111101011110010";
t(525)<="111111111111100011101100";
t(526)<="111111111111011100000000";
t(527)<="111111111111010100111000";
t(528)<="111111111111001110011011";
t(529)<="111111111111001000110000";
t(530)<="111111111111000011111101";
t(531)<="111111111111000000001001";
t(532)<="111111111110111101010111";
t(533)<="111111111110111011101100";
t(534)<="111111111110111011001000";
t(535)<="111111111110111011101110";
t(536)<="111111111110111101011100";
t(537)<="111111111111000000010011";
t(538)<="111111111111000100001110";
t(539)<="111111111111001001001011";
t(540)<="111111111111001111000100";
t(541)<="111111111111010101110011";
t(542)<="111111111111011101010011";
t(543)<="111111111111100101011010";
t(544)<="111111111111101110000001";
t(545)<="111111111111111111111111";
t(546)<="000000000000000000001010";
t(547)<="000000000000001001011000";
t(548)<="000000000000010010100000";
t(549)<="000000000000011011011000";
t(550)<="000000000000100011110111";
t(551)<="000000000000101011110010";
t(552)<="000000000000110011000010";
t(553)<="000000000000111001011111";
t(554)<="000000000000111111000000";
t(555)<="000000000001000011100001";
t(556)<="000000000001000110111100";
t(557)<="000000000001001001001100";
t(558)<="000000000001001010001111";
t(559)<="000000000001001010000011";
t(560)<="000000000001001000101000";
t(561)<="000000000001000101111111";
t(562)<="000000000001000010001011";
t(563)<="000000000000111101001110";
t(564)<="000000000000110111001101";
t(565)<="000000000000110000010000";
t(566)<="000000000000101000011100";
t(567)<="000000000000011111111001";
t(568)<="000000000000010110110001";
t(569)<="000000000000001101001101";
t(570)<="000000000000000011010111";
t(571)<="111111111111111111111111";
t(572)<="111111111111101111011110";
t(573)<="111111111111100101110000";
t(574)<="111111111111011100011011";
t(575)<="111111111111010011101000";
t(576)<="111111111111001011100000";
t(577)<="111111111111000100001101";
t(578)<="111111111110111101110110";
t(579)<="111111111110111000100100";
t(580)<="111111111110110100011100";
t(581)<="111111111110110001100010";
t(582)<="111111111110101111111011";
t(583)<="111111111110101111101001";
t(584)<="111111111110110000101101";
t(585)<="111111111110110011000101";
t(586)<="111111111110110110110001";
t(587)<="111111111110111011101100";
t(588)<="111111111111000001110010";
t(589)<="111111111111001000111110";
t(590)<="111111111111010001000111";
t(591)<="111111111111011010000101";
t(592)<="111111111111100011110000";
t(593)<="111111111111101101111101";
t(594)<="111111111111111111111111";
t(595)<="000000000000000011010011";
t(596)<="000000000000001110000101";
t(597)<="000000000000011000101101";
t(598)<="000000000000100010111111";
t(599)<="000000000000101100110000";
t(600)<="000000000000110101110101";
t(601)<="000000000000111110000101";
t(602)<="000000000001000101010110";
t(603)<="000000000001001011100000";
t(604)<="000000000001010000011100";
t(605)<="000000000001010100000101";
t(606)<="000000000001010110010101";
t(607)<="000000000001010111001010";
t(608)<="000000000001010110100010";
t(609)<="000000000001010100011110";
t(610)<="000000000001010000111111";
t(611)<="000000000001001100000111";
t(612)<="000000000001000101111100";
t(613)<="000000000000111110100100";
t(614)<="000000000000110110000110";
t(615)<="000000000000101100101010";
t(616)<="000000000000100010011011";
t(617)<="000000000000010111100010";
t(618)<="000000000000001100001011";
t(619)<="000000000000000000100011";
t(620)<="111111111111111111111111";
t(621)<="111111111111101001001101";
t(622)<="111111111111011101111001";
t(623)<="111111111111010011000100";
t(624)<="111111111111001000111010";
t(625)<="111111111110111111100111";
t(626)<="111111111110110111010100";
t(627)<="111111111110110000001100";
t(628)<="111111111110101010010101";
t(629)<="111111111110100101110111";
t(630)<="111111111110100010111000";
t(631)<="111111111110100001011010";
t(632)<="111111111110100001100001";
t(633)<="111111111110100011001101";
t(634)<="111111111110100110011101";
t(635)<="111111111110101011001101";
t(636)<="111111111110110001011011";
t(637)<="111111111110111000111111";
t(638)<="111111111111000001110011";
t(639)<="111111111111001011101100";
t(640)<="111111111111010110100011";
t(641)<="111111111111100010001010";
t(642)<="111111111111101110010110";
t(643)<="111111111111111111111111";
t(644)<="000000000000000111101011";
t(645)<="000000000000010100011001";
t(646)<="000000000000100000110110";
t(647)<="000000000000101100110110";
t(648)<="000000000000111000001100";
t(649)<="000000000001000010101011";
t(650)<="000000000001001100001000";
t(651)<="000000000001010100010111";
t(652)<="000000000001011011010000";
t(653)<="000000000001100000101011";
t(654)<="000000000001100100100001";
t(655)<="000000000001100110101110";
t(656)<="000000000001100111001101";
t(657)<="000000000001100101111111";
t(658)<="000000000001100011000011";
t(659)<="000000000001011110011100";
t(660)<="000000000001011000001110";
t(661)<="000000000001010000011111";
t(662)<="000000000001000111010110";
t(663)<="000000000000111100111101";
t(664)<="000000000000110001011110";
t(665)<="000000000000100101000100";
t(666)<="000000000000010111111101";
t(667)<="000000000000001010010110";
t(668)<="111111111111111111111111";
t(669)<="111111111111101110100011";
t(670)<="111111111111100000110100";
t(671)<="111111111111010011011111";
t(672)<="111111111111000110110100";
t(673)<="111111111110111011000000";
t(674)<="111111111110110000010000";
t(675)<="111111111110100110110000";
t(676)<="111111111110011110101011";
t(677)<="111111111110011000001010";
t(678)<="111111111110010011010101";
t(679)<="111111111110010000010001";
t(680)<="111111111110001111000100";
t(681)<="111111111110001111101110";
t(682)<="111111111110010010010001";
t(683)<="111111111110010110101010";
t(684)<="111111111110011100110110";
t(685)<="111111111110100100101111";
t(686)<="111111111110101110001101";
t(687)<="111111111110111001001000";
t(688)<="111111111111000101010011";
t(689)<="111111111111010010100011";
t(690)<="111111111111100000101011";
t(691)<="111111111111101111011010";
t(692)<="111111111111111111111111";
t(693)<="000000000000001101110101";
t(694)<="000000000000011100111111";
t(695)<="000000000000101011110010";
t(696)<="000000000000111001111110";
t(697)<="000000000001000111010011";
t(698)<="000000000001010011100011";
t(699)<="000000000001011110011111";
t(700)<="000000000001100111111100";
t(701)<="000000000001101111101110";
t(702)<="000000000001110101101101";
t(703)<="000000000001111001110010";
t(704)<="000000000001111011110110";
t(705)<="000000000001111011110111";
t(706)<="000000000001111001110011";
t(707)<="000000000001110101101101";
t(708)<="000000000001101111100110";
t(709)<="000000000001100111100110";
t(710)<="000000000001011101110010";
t(711)<="000000000001010010010101";
t(712)<="000000000001000101011010";
t(713)<="000000000000110111001111";
t(714)<="000000000000101000000001";
t(715)<="000000000000011000000000";
t(716)<="000000000000000111011110";
t(717)<="111111111111111111111111";
t(718)<="111111111111100101111001";
t(719)<="111111111111010101011010";
t(720)<="111111111111000101100000";
t(721)<="111111111110110110011101";
t(722)<="111111111110101000100000";
t(723)<="111111111110011011111001";
t(724)<="111111111110010000110111";
t(725)<="111111111110000111100110";
t(726)<="111111111110000000010000";
t(727)<="111111111101111010111111";
t(728)<="111111111101110111111010";
t(729)<="111111111101110111000101";
t(730)<="111111111101111000100001";
t(731)<="111111111101111100001111";
t(732)<="111111111110000010001101";
t(733)<="111111111110001010010100";
t(734)<="111111111110010100011101";
t(735)<="111111111110100000011111";
t(736)<="111111111110101110001101";
t(737)<="111111111110111101011011";
t(738)<="111111111111001101111000";
t(739)<="111111111111011111010100";
t(740)<="111111111111110001011100";
t(741)<="000000000000000011111110";
t(742)<="000000000000010110100111";
t(743)<="000000000000101001000001";
t(744)<="000000000000111010111010";
t(745)<="000000000001001011111110";
t(746)<="000000000001011011111010";
t(747)<="000000000001101010011101";
t(748)<="000000000001110111010111";
t(749)<="000000000010000010011000";
t(750)<="000000000010001011010100";
t(751)<="000000000010010010000000";
t(752)<="000000000010010110010100";
t(753)<="000000000010011000001001";
t(754)<="000000000010010111011101";
t(755)<="000000000010010100001111";
t(756)<="000000000010001110100000";
t(757)<="000000000010000110010110";
t(758)<="000000000001111011110111";
t(759)<="000000000001101111001101";
t(760)<="000000000001100000100110";
t(761)<="000000000001010000001110";
t(762)<="000000000000111110010111";
t(763)<="000000000000101011010011";
t(764)<="000000000000010111010101";
t(765)<="000000000000000010110011";
t(766)<="111111111111101110000001";
t(767)<="111111111111011001010111";
t(768)<="111111111111000101001001";
t(769)<="111111111110110001101110";
t(770)<="111111111110011111011100";
t(771)<="111111111110001110100110";
t(772)<="111111111101111111011111";
t(773)<="111111111101110010011000";
t(774)<="111111111101100111100001";
t(775)<="111111111101011111000111";
t(776)<="111111111101011001010100";
t(777)<="111111111101010110010000";
t(778)<="111111111101010101111111";
t(779)<="111111111101011000100101";
t(780)<="111111111101011101111111";
t(781)<="111111111101100110001011";
t(782)<="111111111101110001000000";
t(783)<="111111111101111110010101";
t(784)<="111111111110001101111110";
t(785)<="111111111110011111101011";
t(786)<="111111111110110011001010";
t(787)<="111111111111001000001000";
t(788)<="111111111111011110010000";
t(789)<="111111111111111111111111";
t(790)<="000000000000001100011111";
t(791)<="000000000000100011110101";
t(792)<="000000000000111010110101";
t(793)<="000000000001010001000100";
t(794)<="000000000001100110001100";
t(795)<="000000000001111001110100";
t(796)<="000000000010001011100111";
t(797)<="000000000010011011010000";
t(798)<="000000000010101000011110";
t(799)<="000000000010110011000000";
t(800)<="000000000010111010101010";
t(801)<="000000000010111111010001";
t(802)<="000000000011000000101110";
t(803)<="000000000010111110111111";
t(804)<="000000000010111010000001";
t(805)<="000000000010110001111001";
t(806)<="000000000010100110101101";
t(807)<="000000000010011000100110";
t(808)<="000000000010000111110011";
t(809)<="000000000001110100100010";
t(810)<="000000000001011111000111";
t(811)<="000000000001000111110111";
t(812)<="000000000000101111001010";
t(813)<="000000000000010101011001";
t(814)<="111111111111111111111111";
t(815)<="111111111111100000010110";
t(816)<="111111111111000101111101";
t(817)<="111111111110101100001111";
t(818)<="111111111110010011101000";
t(819)<="111111111101111100100011";
t(820)<="111111111101100111011010";
t(821)<="111111111101010100100101";
t(822)<="111111111101000100011010";
t(823)<="111111111100110111001011";
t(824)<="111111111100101101001010";
t(825)<="111111111100100110100100";
t(826)<="111111111100100011100001";
t(827)<="111111111100100100001001";
t(828)<="111111111100101000011100";
t(829)<="111111111100110000011010";
t(830)<="111111111100111011111101";
t(831)<="111111111101001010111010";
t(832)<="111111111101011101000101";
t(833)<="111111111101110010001101";
t(834)<="111111111110001001111101";
t(835)<="111111111110100011111111";
t(836)<="111111111110111111111000";
t(837)<="111111111111011101001011";
t(838)<="111111111111111111111111";
t(839)<="000000000000011010001001";
t(840)<="000000000000111000110100";
t(841)<="000000000001010110111010";
t(842)<="000000000001110011111100";
t(843)<="000000000010001111011001";
t(844)<="000000000010101000110011";
t(845)<="000000000010111111101101";
t(846)<="000000000011010011101101";
t(847)<="000000000011100100011011";
t(848)<="000000000011110001100001";
t(849)<="000000000011111010110000";
t(850)<="000000000011111111111001";
t(851)<="000000000100000000110101";
t(852)<="000000000011111101011101";
t(853)<="000000000011110101110011";
t(854)<="000000000011101001111011";
t(855)<="000000000011011001111101";
t(856)<="000000000011000110000111";
t(857)<="000000000010101110101011";
t(858)<="000000000010010011111111";
t(859)<="000000000001110110011100";
t(860)<="000000000001010110011111";
t(861)<="000000000000110100101000";
t(862)<="000000000000010001011001";
t(863)<="111111111111101101011000";
t(864)<="111111111111001001001001";
t(865)<="111111111110100101010010";
t(866)<="111111111110000010011100";
t(867)<="111111111101100001001011";
t(868)<="111111111101000010000101";
t(869)<="111111111100100101101101";
t(870)<="111111111100001100100100";
t(871)<="111111111011110111001000";
t(872)<="111111111011100101110011";
t(873)<="111111111011011000111100";
t(874)<="111111111011010000110101";
t(875)<="111111111011001101101011";
t(876)<="111111111011001111100111";
t(877)<="111111111011010110101100";
t(878)<="111111111011100010110111";
t(879)<="111111111011110100000000";
t(880)<="111111111100001001111100";
t(881)<="111111111100100100010110";
t(882)<="111111111101000010111000";
t(883)<="111111111101100101000101";
t(884)<="111111111110001010011100";
t(885)<="111111111110110010011011";
t(886)<="111111111111011100010111";
t(887)<="000000000000000111101000";
t(888)<="000000000000110011011111";
t(889)<="000000000001011111010000";
t(890)<="000000000010001010001011";
t(891)<="000000000010110011100010";
t(892)<="000000000011011010100110";
t(893)<="000000000011111110101101";
t(894)<="000000000100011111001010";
t(895)<="000000000100111011011001";
t(896)<="000000000101010010110110";
t(897)<="000000000101100101000010";
t(898)<="000000000101110001100011";
t(899)<="000000000101111000000110";
t(900)<="000000000101111000011101";
t(901)<="000000000101110010011111";
t(902)<="000000000101100110001011";
t(903)<="000000000101010011100111";
t(904)<="000000000100111010111110";
t(905)<="000000000100011100100011";
t(906)<="000000000011111000101110";
t(907)<="000000000011010000000000";
t(908)<="000000000010100010111101";
t(909)<="000000000001110010010000";
t(910)<="000000000000111110100111";
t(911)<="000000000000001000110101";
t(912)<="111111111111010001110001";
t(913)<="111111111110011010010011";
t(914)<="111111111101100011010111";
t(915)<="111111111100101101110110";
t(916)<="111111111011111010101101";
t(917)<="111111111011001010110100";
t(918)<="111111111010011111000100";
t(919)<="111111111001111000010000";
t(920)<="111111111001010111001001";
t(921)<="111111111000111100011011";
t(922)<="111111111000101000101100";
t(923)<="111111111000011100011011";
t(924)<="111111111000011000000001";
t(925)<="111111111000011011101110";
t(926)<="111111111000100111101100";
t(927)<="111111111000111011111010";
t(928)<="111111111001011000010001";
t(929)<="111111111001111100011111";
t(930)<="111111111010101000001011";
t(931)<="111111111011011010110100";
t(932)<="111111111100010011110000";
t(933)<="111111111101010010001100";
t(934)<="111111111110010101010001";
t(935)<="111111111111011011111111";
t(936)<="000000000000100101010010";
t(937)<="000000000001110000000010";
t(938)<="000000000010111011000011";
t(939)<="000000000100000101000100";
t(940)<="000000000101001100111000";
t(941)<="000000000110010001001101";
t(942)<="000000000111010000110100";
t(943)<="000000001000001010100011";
t(944)<="000000001000111101001111";
t(945)<="000000001001100111110110";
t(946)<="000000001010001001011010";
t(947)<="000000001010100001000110";
t(948)<="000000001010101110001011";
t(949)<="000000001010110000000100";
t(950)<="000000001010100110011000";
t(951)<="000000001010010000110110";
t(952)<="000000001001101111011011";
t(953)<="000000001001000010001110";
t(954)<="000000001000001001100011";
t(955)<="000000000111000101111000";
t(956)<="000000000101110111111011";
t(957)<="000000000100100000100010";
t(958)<="000000000011000000110001";
t(959)<="000000000001011001110101";
t(960)<="111111111111101101000110";
t(961)<="111111111101111100000101";
t(962)<="111111111100001000011011";
t(963)<="111111111010010011111000";
t(964)<="111111111000100000010000";
t(965)<="111111110110101111011110";
t(966)<="111111110101000011011101";
t(967)<="111111110011011110001001";
t(968)<="111111110010000001100000";
t(969)<="111111110000101111011011";
t(970)<="111111101111101001101111";
t(971)<="111111101110110010001110";
t(972)<="111111101110001010011111";
t(973)<="111111101101110100000100";
t(974)<="111111101101110000010001";
t(975)<="111111101110000000010001";
t(976)<="111111101110100101000001";
t(977)<="111111101111011111010001";
t(978)<="111111110000101111100001";
t(979)<="111111110010010110000001";
t(980)<="111111110100010010110011";
t(981)<="111111110110100101100110";
t(982)<="111111111001001101111001";
t(983)<="111111111100001010111011";
t(984)<="111111111111011011101010";
t(985)<="000000000010111110110011";
t(986)<="000000000110110010110111";
t(987)<="000000001010110110000011";
t(988)<="000000001111000110011100";
t(989)<="000000010011100001111000";
t(990)<="000000011000000110000011";
t(991)<="000000011100110000011111";
t(992)<="000000100001011110101000";
t(993)<="000000100110001101110011";
t(994)<="000000101010111011010001";
t(995)<="000000101111100100010011";
t(996)<="000000110100000110001000";
t(997)<="000000111000011110000011";
t(998)<="000000111100101001011000";
t(999)<="000001000000100101100101";
t(1000)<="000001000100010000001110";
t(1001)<="000001000111100111000000";
t(1002)<="000001001010100111110101";
t(1003)<="000001001101010000110101";
t(1004)<="000001001111100000010011";
t(1005)<="000001010001010100110100";
t(1006)<="000001010010101101010000";
t(1007)<="000001010011101000101101";
t(1008)<="000001010100000110100100";
t(1009)<="000001010100000110100100";
t(1010)<="000001010011101000101101";
t(1011)<="000001010010101101010000";
t(1012)<="000001010001010100110100";
t(1013)<="000001001111100000010011";
t(1014)<="000001001101010000110101";
t(1015)<="000001001010100111110101";
t(1016)<="000001000111100111000000";
t(1017)<="000001000100010000001110";
t(1018)<="000001000000100101100101";
t(1019)<="000000111100101001011000";
t(1020)<="000000111000011110000011";
t(1021)<="000000110100000110001000";
t(1022)<="000000101111100100010011";
t(1023)<="000000101010111011010001";
t(1024)<="000000100110001101110011";
t(1025)<="000000100001011110101000";
t(1026)<="000000011100110000011111";
t(1027)<="000000011000000110000011";
t(1028)<="000000010011100001111000";
t(1029)<="000000001111000110011100";
t(1030)<="000000001010110110000011";
t(1031)<="000000000110110010110111";
t(1032)<="000000000010111110110011";
t(1033)<="111111111111011011101010";
t(1034)<="111111111100001010111011";
t(1035)<="111111111001001101111001";
t(1036)<="111111110110100101100110";
t(1037)<="111111110100010010110011";
t(1038)<="111111110010010110000001";
t(1039)<="111111110000101111100001";
t(1040)<="111111101111011111010001";
t(1041)<="111111101110100101000001";
t(1042)<="111111101110000000010001";
t(1043)<="111111101101110000010001";
t(1044)<="111111101101110100000100";
t(1045)<="111111101110001010011111";
t(1046)<="111111101110110010001110";
t(1047)<="111111101111101001101111";
t(1048)<="111111110000101111011011";
t(1049)<="111111110010000001100000";
t(1050)<="111111110011011110001001";
t(1051)<="111111110101000011011101";
t(1052)<="111111110110101111011110";
t(1053)<="111111111000100000010000";
t(1054)<="111111111010010011111000";
t(1055)<="111111111100001000011011";
t(1056)<="111111111101111100000101";
t(1057)<="111111111111101101000110";
t(1058)<="000000000001011001110101";
t(1059)<="000000000011000000110001";
t(1060)<="000000000100100000100010";
t(1061)<="000000000101110111111011";
t(1062)<="000000000111000101111000";
t(1063)<="000000001000001001100011";
t(1064)<="000000001001000010001110";
t(1065)<="000000001001101111011011";
t(1066)<="000000001010010000110110";
t(1067)<="000000001010100110011000";
t(1068)<="000000001010110000000100";
t(1069)<="000000001010101110001011";
t(1070)<="000000001010100001000110";
t(1071)<="000000001010001001011010";
t(1072)<="000000001001100111110110";
t(1073)<="000000001000111101001111";
t(1074)<="000000001000001010100011";
t(1075)<="000000000111010000110100";
t(1076)<="000000000110010001001101";
t(1077)<="000000000101001100111000";
t(1078)<="000000000100000101000100";
t(1079)<="000000000010111011000011";
t(1080)<="000000000001110000000010";
t(1081)<="000000000000100101010010";
t(1082)<="111111111111011011111111";
t(1083)<="111111111110010101010001";
t(1084)<="111111111101010010001100";
t(1085)<="111111111100010011110000";
t(1086)<="111111111011011010110100";
t(1087)<="111111111010101000001011";
t(1088)<="111111111001111100011111";
t(1089)<="111111111001011000010001";
t(1090)<="111111111000111011111010";
t(1091)<="111111111000100111101100";
t(1092)<="111111111000011011101110";
t(1093)<="111111111000011000000001";
t(1094)<="111111111000011100011011";
t(1095)<="111111111000101000101100";
t(1096)<="111111111000111100011011";
t(1097)<="111111111001010111001001";
t(1098)<="111111111001111000010000";
t(1099)<="111111111010011111000100";
t(1100)<="111111111011001010110100";
t(1101)<="111111111011111010101101";
t(1102)<="111111111100101101110110";
t(1103)<="111111111101100011010111";
t(1104)<="111111111110011010010011";
t(1105)<="111111111111010001110001";
t(1106)<="000000000000001000110101";
t(1107)<="000000000000111110100111";
t(1108)<="000000000001110010010000";
t(1109)<="000000000010100010111101";
t(1110)<="000000000011010000000000";
t(1111)<="000000000011111000101110";
t(1112)<="000000000100011100100011";
t(1113)<="000000000100111010111110";
t(1114)<="000000000101010011100111";
t(1115)<="000000000101100110001011";
t(1116)<="000000000101110010011111";
t(1117)<="000000000101111000011101";
t(1118)<="000000000101111000000110";
t(1119)<="000000000101110001100011";
t(1120)<="000000000101100101000010";
t(1121)<="000000000101010010110110";
t(1122)<="000000000100111011011001";
t(1123)<="000000000100011111001010";
t(1124)<="000000000011111110101101";
t(1125)<="000000000011011010100110";
t(1126)<="000000000010110011100010";
t(1127)<="000000000010001010001011";
t(1128)<="000000000001011111010000";
t(1129)<="000000000000110011011111";
t(1130)<="000000000000000111101000";
t(1131)<="111111111111011100010111";
t(1132)<="111111111110110010011011";
t(1133)<="111111111110001010011100";
t(1134)<="111111111101100101000101";
t(1135)<="111111111101000010111000";
t(1136)<="111111111100100100010110";
t(1137)<="111111111100001001111100";
t(1138)<="111111111011110100000000";
t(1139)<="111111111011100010110111";
t(1140)<="111111111011010110101100";
t(1141)<="111111111011001111100111";
t(1142)<="111111111011001101101011";
t(1143)<="111111111011010000110101";
t(1144)<="111111111011011000111100";
t(1145)<="111111111011100101110011";
t(1146)<="111111111011110111001000";
t(1147)<="111111111100001100100100";
t(1148)<="111111111100100101101101";
t(1149)<="111111111101000010000101";
t(1150)<="111111111101100001001011";
t(1151)<="111111111110000010011100";
t(1152)<="111111111110100101010010";
t(1153)<="111111111111001001001001";
t(1154)<="111111111111101101011000";
t(1155)<="000000000000010001011001";
t(1156)<="000000000000110100101000";
t(1157)<="000000000001010110011111";
t(1158)<="000000000001110110011100";
t(1159)<="000000000010010011111111";
t(1160)<="000000000010101110101011";
t(1161)<="000000000011000110000111";
t(1162)<="000000000011011001111101";
t(1163)<="000000000011101001111011";
t(1164)<="000000000011110101110011";
t(1165)<="000000000011111101011101";
t(1166)<="000000000100000000110101";
t(1167)<="000000000011111111111001";
t(1168)<="000000000011111010110000";
t(1169)<="000000000011110001100001";
t(1170)<="000000000011100100011011";
t(1171)<="000000000011010011101101";
t(1172)<="000000000010111111101101";
t(1173)<="000000000010101000110011";
t(1174)<="000000000010001111011001";
t(1175)<="000000000001110011111100";
t(1176)<="000000000001010110111010";
t(1177)<="000000000000111000110100";
t(1178)<="000000000000011010001001";
t(1179)<="111111111111111111111111";
t(1180)<="111111111111011101001011";
t(1181)<="111111111110111111111000";
t(1182)<="111111111110100011111111";
t(1183)<="111111111110001001111101";
t(1184)<="111111111101110010001101";
t(1185)<="111111111101011101000101";
t(1186)<="111111111101001010111010";
t(1187)<="111111111100111011111101";
t(1188)<="111111111100110000011010";
t(1189)<="111111111100101000011100";
t(1190)<="111111111100100100001001";
t(1191)<="111111111100100011100001";
t(1192)<="111111111100100110100100";
t(1193)<="111111111100101101001010";
t(1194)<="111111111100110111001011";
t(1195)<="111111111101000100011010";
t(1196)<="111111111101010100100101";
t(1197)<="111111111101100111011010";
t(1198)<="111111111101111100100011";
t(1199)<="111111111110010011101000";
t(1200)<="111111111110101100001111";
t(1201)<="111111111111000101111101";
t(1202)<="111111111111100000010110";
t(1203)<="111111111111111111111111";
t(1204)<="000000000000010101011001";
t(1205)<="000000000000101111001010";
t(1206)<="000000000001000111110111";
t(1207)<="000000000001011111000111";
t(1208)<="000000000001110100100010";
t(1209)<="000000000010000111110011";
t(1210)<="000000000010011000100110";
t(1211)<="000000000010100110101101";
t(1212)<="000000000010110001111001";
t(1213)<="000000000010111010000001";
t(1214)<="000000000010111110111111";
t(1215)<="000000000011000000101110";
t(1216)<="000000000010111111010001";
t(1217)<="000000000010111010101010";
t(1218)<="000000000010110011000000";
t(1219)<="000000000010101000011110";
t(1220)<="000000000010011011010000";
t(1221)<="000000000010001011100111";
t(1222)<="000000000001111001110100";
t(1223)<="000000000001100110001100";
t(1224)<="000000000001010001000100";
t(1225)<="000000000000111010110101";
t(1226)<="000000000000100011110101";
t(1227)<="000000000000001100011111";
t(1228)<="111111111111111111111111";
t(1229)<="111111111111011110010000";
t(1230)<="111111111111001000001000";
t(1231)<="111111111110110011001010";
t(1232)<="111111111110011111101011";
t(1233)<="111111111110001101111110";
t(1234)<="111111111101111110010101";
t(1235)<="111111111101110001000000";
t(1236)<="111111111101100110001011";
t(1237)<="111111111101011101111111";
t(1238)<="111111111101011000100101";
t(1239)<="111111111101010101111111";
t(1240)<="111111111101010110010000";
t(1241)<="111111111101011001010100";
t(1242)<="111111111101011111000111";
t(1243)<="111111111101100111100001";
t(1244)<="111111111101110010011000";
t(1245)<="111111111101111111011111";
t(1246)<="111111111110001110100110";
t(1247)<="111111111110011111011100";
t(1248)<="111111111110110001101110";
t(1249)<="111111111111000101001001";
t(1250)<="111111111111011001010111";
t(1251)<="111111111111101110000001";
t(1252)<="000000000000000010110011";
t(1253)<="000000000000010111010101";
t(1254)<="000000000000101011010011";
t(1255)<="000000000000111110010111";
t(1256)<="000000000001010000001110";
t(1257)<="000000000001100000100110";
t(1258)<="000000000001101111001101";
t(1259)<="000000000001111011110111";
t(1260)<="000000000010000110010110";
t(1261)<="000000000010001110100000";
t(1262)<="000000000010010100001111";
t(1263)<="000000000010010111011101";
t(1264)<="000000000010011000001001";
t(1265)<="000000000010010110010100";
t(1266)<="000000000010010010000000";
t(1267)<="000000000010001011010100";
t(1268)<="000000000010000010011000";
t(1269)<="000000000001110111010111";
t(1270)<="000000000001101010011101";
t(1271)<="000000000001011011111010";
t(1272)<="000000000001001011111110";
t(1273)<="000000000000111010111010";
t(1274)<="000000000000101001000001";
t(1275)<="000000000000010110100111";
t(1276)<="000000000000000011111110";
t(1277)<="111111111111110001011100";
t(1278)<="111111111111011111010100";
t(1279)<="111111111111001101111000";
t(1280)<="111111111110111101011011";
t(1281)<="111111111110101110001101";
t(1282)<="111111111110100000011111";
t(1283)<="111111111110010100011101";
t(1284)<="111111111110001010010100";
t(1285)<="111111111110000010001101";
t(1286)<="111111111101111100001111";
t(1287)<="111111111101111000100001";
t(1288)<="111111111101110111000101";
t(1289)<="111111111101110111111010";
t(1290)<="111111111101111010111111";
t(1291)<="111111111110000000010000";
t(1292)<="111111111110000111100110";
t(1293)<="111111111110010000110111";
t(1294)<="111111111110011011111001";
t(1295)<="111111111110101000100000";
t(1296)<="111111111110110110011101";
t(1297)<="111111111111000101100000";
t(1298)<="111111111111010101011010";
t(1299)<="111111111111100101111001";
t(1300)<="111111111111111111111111";
t(1301)<="000000000000000111011110";
t(1302)<="000000000000011000000000";
t(1303)<="000000000000101000000001";
t(1304)<="000000000000110111001111";
t(1305)<="000000000001000101011010";
t(1306)<="000000000001010010010101";
t(1307)<="000000000001011101110010";
t(1308)<="000000000001100111100110";
t(1309)<="000000000001101111100110";
t(1310)<="000000000001110101101101";
t(1311)<="000000000001111001110011";
t(1312)<="000000000001111011110111";
t(1313)<="000000000001111011110110";
t(1314)<="000000000001111001110010";
t(1315)<="000000000001110101101101";
t(1316)<="000000000001101111101110";
t(1317)<="000000000001100111111100";
t(1318)<="000000000001011110011111";
t(1319)<="000000000001010011100011";
t(1320)<="000000000001000111010011";
t(1321)<="000000000000111001111110";
t(1322)<="000000000000101011110010";
t(1323)<="000000000000011100111111";
t(1324)<="000000000000001101110101";
t(1325)<="111111111111111111111111";
t(1326)<="111111111111101111011010";
t(1327)<="111111111111100000101011";
t(1328)<="111111111111010010100011";
t(1329)<="111111111111000101010011";
t(1330)<="111111111110111001001000";
t(1331)<="111111111110101110001101";
t(1332)<="111111111110100100101111";
t(1333)<="111111111110011100110110";
t(1334)<="111111111110010110101010";
t(1335)<="111111111110010010010001";
t(1336)<="111111111110001111101110";
t(1337)<="111111111110001111000100";
t(1338)<="111111111110010000010001";
t(1339)<="111111111110010011010101";
t(1340)<="111111111110011000001010";
t(1341)<="111111111110011110101011";
t(1342)<="111111111110100110110000";
t(1343)<="111111111110110000010000";
t(1344)<="111111111110111011000000";
t(1345)<="111111111111000110110100";
t(1346)<="111111111111010011011111";
t(1347)<="111111111111100000110100";
t(1348)<="111111111111101110100011";
t(1349)<="111111111111111111111111";
t(1350)<="000000000000001010010110";
t(1351)<="000000000000010111111101";
t(1352)<="000000000000100101000100";
t(1353)<="000000000000110001011110";
t(1354)<="000000000000111100111101";
t(1355)<="000000000001000111010110";
t(1356)<="000000000001010000011111";
t(1357)<="000000000001011000001110";
t(1358)<="000000000001011110011100";
t(1359)<="000000000001100011000011";
t(1360)<="000000000001100101111111";
t(1361)<="000000000001100111001101";
t(1362)<="000000000001100110101110";
t(1363)<="000000000001100100100001";
t(1364)<="000000000001100000101011";
t(1365)<="000000000001011011010000";
t(1366)<="000000000001010100010111";
t(1367)<="000000000001001100001000";
t(1368)<="000000000001000010101011";
t(1369)<="000000000000111000001100";
t(1370)<="000000000000101100110110";
t(1371)<="000000000000100000110110";
t(1372)<="000000000000010100011001";
t(1373)<="000000000000000111101011";
t(1374)<="111111111111111111111111";
t(1375)<="111111111111101110010110";
t(1376)<="111111111111100010001010";
t(1377)<="111111111111010110100011";
t(1378)<="111111111111001011101100";
t(1379)<="111111111111000001110011";
t(1380)<="111111111110111000111111";
t(1381)<="111111111110110001011011";
t(1382)<="111111111110101011001101";
t(1383)<="111111111110100110011101";
t(1384)<="111111111110100011001101";
t(1385)<="111111111110100001100001";
t(1386)<="111111111110100001011010";
t(1387)<="111111111110100010111000";
t(1388)<="111111111110100101110111";
t(1389)<="111111111110101010010101";
t(1390)<="111111111110110000001100";
t(1391)<="111111111110110111010100";
t(1392)<="111111111110111111100111";
t(1393)<="111111111111001000111010";
t(1394)<="111111111111010011000100";
t(1395)<="111111111111011101111001";
t(1396)<="111111111111101001001101";
t(1397)<="111111111111111111111111";
t(1398)<="000000000000000000100011";
t(1399)<="000000000000001100001011";
t(1400)<="000000000000010111100010";
t(1401)<="000000000000100010011011";
t(1402)<="000000000000101100101010";
t(1403)<="000000000000110110000110";
t(1404)<="000000000000111110100100";
t(1405)<="000000000001000101111100";
t(1406)<="000000000001001100000111";
t(1407)<="000000000001010000111111";
t(1408)<="000000000001010100011110";
t(1409)<="000000000001010110100010";
t(1410)<="000000000001010111001010";
t(1411)<="000000000001010110010101";
t(1412)<="000000000001010100000101";
t(1413)<="000000000001010000011100";
t(1414)<="000000000001001011100000";
t(1415)<="000000000001000101010110";
t(1416)<="000000000000111110000101";
t(1417)<="000000000000110101110101";
t(1418)<="000000000000101100110000";
t(1419)<="000000000000100010111111";
t(1420)<="000000000000011000101101";
t(1421)<="000000000000001110000101";
t(1422)<="000000000000000011010011";
t(1423)<="111111111111111111111111";
t(1424)<="111111111111101101111101";
t(1425)<="111111111111100011110000";
t(1426)<="111111111111011010000101";
t(1427)<="111111111111010001000111";
t(1428)<="111111111111001000111110";
t(1429)<="111111111111000001110010";
t(1430)<="111111111110111011101100";
t(1431)<="111111111110110110110001";
t(1432)<="111111111110110011000101";
t(1433)<="111111111110110000101101";
t(1434)<="111111111110101111101001";
t(1435)<="111111111110101111111011";
t(1436)<="111111111110110001100010";
t(1437)<="111111111110110100011100";
t(1438)<="111111111110111000100100";
t(1439)<="111111111110111101110110";
t(1440)<="111111111111000100001101";
t(1441)<="111111111111001011100000";
t(1442)<="111111111111010011101000";
t(1443)<="111111111111011100011011";
t(1444)<="111111111111100101110000";
t(1445)<="111111111111101111011110";
t(1446)<="111111111111111111111111";
t(1447)<="000000000000000011010111";
t(1448)<="000000000000001101001101";
t(1449)<="000000000000010110110001";
t(1450)<="000000000000011111111001";
t(1451)<="000000000000101000011100";
t(1452)<="000000000000110000010000";
t(1453)<="000000000000110111001101";
t(1454)<="000000000000111101001110";
t(1455)<="000000000001000010001011";
t(1456)<="000000000001000101111111";
t(1457)<="000000000001001000101000";
t(1458)<="000000000001001010000011";
t(1459)<="000000000001001010001111";
t(1460)<="000000000001001001001100";
t(1461)<="000000000001000110111100";
t(1462)<="000000000001000011100001";
t(1463)<="000000000000111111000000";
t(1464)<="000000000000111001011111";
t(1465)<="000000000000110011000010";
t(1466)<="000000000000101011110010";
t(1467)<="000000000000100011110111";
t(1468)<="000000000000011011011000";
t(1469)<="000000000000010010100000";
t(1470)<="000000000000001001011000";
t(1471)<="000000000000000000001010";
t(1472)<="111111111111111111111111";
t(1473)<="111111111111101110000001";
t(1474)<="111111111111100101011010";
t(1475)<="111111111111011101010011";
t(1476)<="111111111111010101110011";
t(1477)<="111111111111001111000100";
t(1478)<="111111111111001001001011";
t(1479)<="111111111111000100001110";
t(1480)<="111111111111000000010011";
t(1481)<="111111111110111101011100";
t(1482)<="111111111110111011101110";
t(1483)<="111111111110111011001000";
t(1484)<="111111111110111011101100";
t(1485)<="111111111110111101010111";
t(1486)<="111111111111000000001001";
t(1487)<="111111111111000011111101";
t(1488)<="111111111111001000110000";
t(1489)<="111111111111001110011011";
t(1490)<="111111111111010100111000";
t(1491)<="111111111111011100000000";
t(1492)<="111111111111100011101100";
t(1493)<="111111111111101011110010";
t(1494)<="111111111111111111111111";
t(1495)<="111111111111111111111111";
t(1496)<="000000000000000101001111";
t(1497)<="000000000000001101101000";
t(1498)<="000000000000010101110000";
t(1499)<="000000000000011101011101";
t(1500)<="000000000000100100100111";
t(1501)<="000000000000101011001001";
t(1502)<="000000000000110000111001";
t(1503)<="000000000000110101110100";
t(1504)<="000000000000111001110100";
t(1505)<="000000000000111100110101";
t(1506)<="000000000000111110110100";
t(1507)<="000000000000111111110000";
t(1508)<="000000000000111111100111";
t(1509)<="000000000000111110011100";
t(1510)<="000000000000111100001111";
t(1511)<="000000000000111001000010";
t(1512)<="000000000000110100111011";
t(1513)<="000000000000101111111101";
t(1514)<="000000000000101010001110";
t(1515)<="000000000000100011110101";
t(1516)<="000000000000011100111000";
t(1517)<="000000000000010101011111";
t(1518)<="000000000000001101110010";
t(1519)<="000000000000000101111010";
t(1520)<="111111111111111111111111";
t(1521)<="111111111111111111111111";
t(1522)<="111111111111101110011111";
t(1523)<="111111111111100111001011";
t(1524)<="111111111111100000010101";
t(1525)<="111111111111011010000011";
t(1526)<="111111111111010100011011";
t(1527)<="111111111111001111100100";
t(1528)<="111111111111001011100010";
t(1529)<="111111111111001000011001";
t(1530)<="111111111111000110001100";
t(1531)<="111111111111000100111110";
t(1532)<="111111111111000100101110";
t(1533)<="111111111111000101011101";
t(1534)<="111111111111000111001010";
t(1535)<="111111111111001001110010";
t(1536)<="111111111111001101010011";
t(1537)<="111111111111010001101001";
t(1538)<="111111111111010110101101";
t(1539)<="111111111111011100011100";
t(1540)<="111111111111100010101101";
t(1541)<="111111111111101001011100";
t(1542)<="111111111111110000100000";
t(1543)<="111111111111111111111111";
t(1544)<="111111111111111111111111";
t(1545)<="000000000000000110011110";
t(1546)<="000000000000001101101010";
t(1547)<="000000000000010100100100";
t(1548)<="000000000000011011000111";
t(1549)<="000000000000100001001001";
t(1550)<="000000000000100110100111";
t(1551)<="000000000000101011011001";
t(1552)<="000000000000101111011100";
t(1553)<="000000000000110010101011";
t(1554)<="000000000000110101000011";
t(1555)<="000000000000110110100001";
t(1556)<="000000000000110111000110";
t(1557)<="000000000000110110110000";
t(1558)<="000000000000110101100000";
t(1559)<="000000000000110011010111";
t(1560)<="000000000000110000011001";
t(1561)<="000000000000101100101001";
t(1562)<="000000000000101000001011";
t(1563)<="000000000000100011000100";
t(1564)<="000000000000011101011010";
t(1565)<="000000000000010111010011";
t(1566)<="000000000000010000110110";
t(1567)<="000000000000001010001001";
t(1568)<="000000000000000011010100";
t(1569)<="111111111111111111111111";
t(1570)<="111111111111111111111111";
t(1571)<="111111111111101111001011";
t(1572)<="111111111111101000111101";
t(1573)<="111111111111100011001010";
t(1574)<="111111111111011101110111";
t(1575)<="111111111111011001001011";
t(1576)<="111111111111010101001001";
t(1577)<="111111111111010001110111";
t(1578)<="111111111111001111010110";
t(1579)<="111111111111001101101010";
t(1580)<="111111111111001100110100";
t(1581)<="111111111111001100110100";
t(1582)<="111111111111001101101011";
t(1583)<="111111111111001111010111";
t(1584)<="111111111111010001110101";
t(1585)<="111111111111010101000100";
t(1586)<="111111111111011000111111";
t(1587)<="111111111111011101100001";
t(1588)<="111111111111100010100111";
t(1589)<="111111111111101000001010";
t(1590)<="111111111111101110000100";
t(1591)<="111111111111111111111111";
t(1592)<="111111111111111111111111";
t(1593)<="000000000000000000111100";
t(1594)<="000000000000000111010001";
t(1595)<="000000000000001101011100";
t(1596)<="000000000000010011010110";
t(1597)<="000000000000011000111010";
t(1598)<="000000000000011110000001";
t(1599)<="000000000000100010100111";
t(1600)<="000000000000100110100110";
t(1601)<="000000000000101001111011";
t(1602)<="000000000000101100100010";
t(1603)<="000000000000101110011001";
t(1604)<="000000000000101111011110";
t(1605)<="000000000000101111110001";
t(1606)<="000000000000101111010001";
t(1607)<="000000000000101101111111";
t(1608)<="000000000000101011111100";
t(1609)<="000000000000101001001100";
t(1610)<="000000000000100101110001";
t(1611)<="000000000000100001110000";
t(1612)<="000000000000011101001100";
t(1613)<="000000000000011000001011";
t(1614)<="000000000000010010110001";
t(1615)<="000000000000001101000111";
t(1616)<="000000000000000111010000";
t(1617)<="000000000000000001010100";
t(1618)<="111111111111111111111111";
t(1619)<="111111111111111111111111";
t(1620)<="111111111111101111111100";
t(1621)<="111111111111101010101000";
t(1622)<="111111111111100101101100";
t(1623)<="111111111111100001001110";
t(1624)<="111111111111011101010010";
t(1625)<="111111111111011001111101";
t(1626)<="111111111111010111010001";
t(1627)<="111111111111010101010001";
t(1628)<="111111111111010011111111";
t(1629)<="111111111111010011011100";
t(1630)<="111111111111010011101001";
t(1631)<="111111111111010100100100";
t(1632)<="111111111111010110001101";
t(1633)<="111111111111011000100010";
t(1634)<="111111111111011011100000";
t(1635)<="111111111111011111000100";
t(1636)<="111111111111100011001001";
t(1637)<="111111111111100111101100";
t(1638)<="111111111111101100100110";
t(1639)<="111111111111110001110100";
t(1640)<="111111111111111111111111";
t(1641)<="111111111111111111111111";
t(1642)<="000000000000000010010100";
t(1643)<="000000000000000111110011";
t(1644)<="000000000000001101001000";
t(1645)<="000000000000010010001101";
t(1646)<="000000000000010110111101";
t(1647)<="000000000000011011010011";
t(1648)<="000000000000011111001011";
t(1649)<="000000000000100010100000";
t(1650)<="000000000000100101010000";
t(1651)<="000000000000100111010111";
t(1652)<="000000000000101000110100";
t(1653)<="000000000000101001100101";
t(1654)<="000000000000101001101001";
t(1655)<="000000000000101001000010";
t(1656)<="000000000000100111101111";
t(1657)<="000000000000100101110011";
t(1658)<="000000000000100011001111";
t(1659)<="000000000000100000000110";
t(1660)<="000000000000011100011101";
t(1661)<="000000000000011000010111";
t(1662)<="000000000000010011111000";
t(1663)<="000000000000001111000110";
t(1664)<="000000000000001010000101";
t(1665)<="000000000000000100111100";
t(1666)<="111111111111111111111111";
t(1667)<="111111111111111111111111";
t(1668)<="111111111111111111111111";
t(1669)<="111111111111110000101001";
t(1670)<="111111111111101100000101";
t(1671)<="111111111111100111110110";
t(1672)<="111111111111100100000011";
t(1673)<="111111111111100000101111";
t(1674)<="111111111111011101111100";
t(1675)<="111111111111011011101111";
t(1676)<="111111111111011010001001";
t(1677)<="111111111111011001001100";
t(1678)<="111111111111011000111000";
t(1679)<="111111111111011001001101";
t(1680)<="111111111111011010001100";
t(1681)<="111111111111011011110010";
t(1682)<="111111111111011101111110";
t(1683)<="111111111111100000101101";
t(1684)<="111111111111100011111101";
t(1685)<="111111111111100111101001";
t(1686)<="111111111111101011101110";
t(1687)<="111111111111110000000111";
t(1688)<="111111111111111111111111";
t(1689)<="111111111111111111111111";
t(1690)<="111111111111111111111111";
t(1691)<="000000000000000011010010";
t(1692)<="000000000000001000000101";
t(1693)<="000000000000001100101111";
t(1694)<="000000000000010001001000";
t(1695)<="000000000000010101001111";
t(1696)<="000000000000011000111110";
t(1697)<="000000000000011100010001";
t(1698)<="000000000000011111000101";
t(1699)<="000000000000100001010111";
t(1700)<="000000000000100011000101";
t(1701)<="000000000000100100001101";
t(1702)<="000000000000100100101111";
t(1703)<="000000000000100100101010";
t(1704)<="000000000000100011111101";
t(1705)<="000000000000100010101011";
t(1706)<="000000000000100000110101";
t(1707)<="000000000000011110011100";
t(1708)<="000000000000011011100100";
t(1709)<="000000000000011000001111";
t(1710)<="000000000000010100100010";
t(1711)<="000000000000010000100000";
t(1712)<="000000000000001100001110";
t(1713)<="000000000000000111110000";
t(1714)<="000000000000000011001011";
t(1715)<="111111111111111111111111";
t(1716)<="111111111111111111111111";
t(1717)<="111111111111111111111111";
t(1718)<="111111111111110001010101";
t(1719)<="111111111111101101010110";
t(1720)<="111111111111101001101100";
t(1721)<="111111111111100110011011";
t(1722)<="111111111111100011100110";
t(1723)<="111111111111100001010000";
t(1724)<="111111111111011111011011";
t(1725)<="111111111111011110001001";
t(1726)<="111111111111011101011011";
t(1727)<="111111111111011101010011";
t(1728)<="111111111111011101101111";
t(1729)<="111111111111011110101111";
t(1730)<="111111111111100000010010";
t(1731)<="111111111111100010010111";
t(1732)<="111111111111100100111010";
t(1733)<="111111111111100111111001";
t(1734)<="111111111111101011010001";
t(1735)<="111111111111101110111110";
t(1736)<="111111111111111111111111";
t(1737)<="111111111111111111111111";
t(1738)<="111111111111111111111111";
t(1739)<="111111111111111111111111";
t(1740)<="000000000000000100001000";
t(1741)<="000000000000001000011000";
t(1742)<="000000000000001100011111";
t(1743)<="000000000000010000010111";
t(1744)<="000000000000010011111101";
t(1745)<="000000000000010111001101";
t(1746)<="000000000000011010000011";
t(1747)<="000000000000011100011110";
t(1748)<="000000000000011110011001";
t(1749)<="000000000000011111110100";
t(1750)<="000000000000100000101100";
t(1751)<="000000000000100001000010";
t(1752)<="000000000000100000110101";
t(1753)<="000000000000100000000101";
t(1754)<="000000000000011110110011";
t(1755)<="000000000000011101000001";
t(1756)<="000000000000011010110001";
t(1757)<="000000000000011000000100";
t(1758)<="000000000000010100111111";
t(1759)<="000000000000010001100101";
t(1760)<="000000000000001101111000";
t(1761)<="000000000000001001111110";
t(1762)<="000000000000000101111010";
t(1763)<="000000000000000001110001";
t(1764)<="111111111111111111111111";
t(1765)<="111111111111111111111111";
t(1766)<="111111111111111111111111";
t(1767)<="111111111111110001101101";
t(1768)<="111111111111101110001010";
t(1769)<="111111111111101010111011";
t(1770)<="111111111111101000000010";
t(1771)<="111111111111100101100100";
t(1772)<="111111111111100011100010";
t(1773)<="111111111111100001111110";
t(1774)<="111111111111100000111011";
t(1775)<="111111111111100000011001";
t(1776)<="111111111111100000011000";
t(1777)<="111111111111100000111001";
t(1778)<="111111111111100001111011";
t(1779)<="111111111111100011011100";
t(1780)<="111111111111100101011011";
t(1781)<="111111111111100111110111";
t(1782)<="111111111111101010101011";
t(1783)<="111111111111101101110101";
t(1784)<="111111111111110001010010";
t(1785)<="111111111111111111111111";
t(1786)<="111111111111111111111111";
t(1787)<="111111111111111111111111";
t(1788)<="000000000000000000110101";
t(1789)<="000000000000000100110100";
t(1790)<="000000000000001000101110";
t(1791)<="000000000000001100011110";
t(1792)<="000000000000010000000000";
t(1793)<="000000000000010011010001";
t(1794)<="000000000000010110001100";
t(1795)<="000000000000011000110001";
t(1796)<="000000000000011010111010";
t(1797)<="000000000000011100100111";
t(1798)<="000000000000011101110101";
t(1799)<="000000000000011110100100";
t(1800)<="000000000000011110110010";
t(1801)<="000000000000011110100000";
t(1802)<="000000000000011101101101";
t(1803)<="000000000000011100011100";
t(1804)<="000000000000011010101100";
t(1805)<="000000000000011000100000";
t(1806)<="000000000000010101111010";
t(1807)<="000000000000010010111110";
t(1808)<="000000000000001111101101";
t(1809)<="000000000000001100001101";
t(1810)<="000000000000001000011111";
t(1811)<="000000000000000100101001";
t(1812)<="000000000000000000101110";
t(1813)<="111111111111111111111111";
t(1814)<="111111111111111111111111";
t(1815)<="111111111111111111111111";
t(1816)<="111111111111110001100110";
t(1817)<="111111111111101110010001";
t(1818)<="111111111111101011001111";
t(1819)<="111111111111101000100010";
t(1820)<="111111111111100110001111";
t(1821)<="111111111111100100010110";
t(1822)<="111111111111100010111011";
t(1823)<="111111111111100001111110";
t(1824)<="111111111111100001100001";
t(1825)<="111111111111100001100100";
t(1826)<="111111111111100010000111";
t(1827)<="111111111111100011001010";
t(1828)<="111111111111100100101011";
t(1829)<="111111111111100110101001";
t(1830)<="111111111111101001000001";
t(1831)<="111111111111101011110010";
t(1832)<="111111111111101110111000";
t(1833)<="111111111111110010010000";
t(1834)<="111111111111111111111111";
t(1835)<="111111111111111111111111";
t(1836)<="111111111111111111111111";
t(1837)<="000000000000000001011101";
t(1838)<="000000000000000101010111";
t(1839)<="000000000000001001001101";
t(1840)<="000000000000001100111000";
t(1841)<="000000000000010000010111";
t(1842)<="000000000000010011100101";
t(1843)<="000000000000010110011111";
t(1844)<="000000000000011001000001";
t(1845)<="000000000000011011001010";
t(1846)<="000000000000011100110111";
t(1847)<="000000000000011110000101";
t(1848)<="000000000000011110110101";
t(1849)<="000000000000011111000100";
t(1850)<="000000000000011110110011";
t(1851)<="000000000000011110000010";
t(1852)<="000000000000011100110001";
t(1853)<="000000000000011011000010";
t(1854)<="000000000000011000110111";
t(1855)<="000000000000010110010001";
t(1856)<="000000000000010011010011";
t(1857)<="000000000000010000000001";
t(1858)<="000000000000001100011101";
t(1859)<="000000000000001000101100";
t(1860)<="000000000000000100110000";
t(1861)<="000000000000000000101111";
t(1862)<="111111111111111111111111";
t(1863)<="111111111111111111111111";
t(1864)<="111111111111111111111111";
t(1865)<="111111111111110001000001";
t(1866)<="111111111111101101011111";
t(1867)<="111111111111101010010000";
t(1868)<="111111111111100111010110";
t(1869)<="111111111111100100110100";
t(1870)<="111111111111100010101110";
t(1871)<="111111111111100001000101";
t(1872)<="111111111111011111111011";
t(1873)<="111111111111011111010011";
t(1874)<="111111111111011111001011";
t(1875)<="111111111111011111100101";
t(1876)<="111111111111100000100000";
t(1877)<="111111111111100001111101";
t(1878)<="111111111111100011111000";
t(1879)<="111111111111100110010001";
t(1880)<="111111111111101001000110";
t(1881)<="111111111111101100010011";
t(1882)<="111111111111101111110110";
t(1883)<="111111111111111111111111";
t(1884)<="111111111111111111111111";
t(1885)<="111111111111111111111111";
t(1886)<="000000000000000000010000";
t(1887)<="000000000000000100100110";
t(1888)<="000000000000001000111001";
t(1889)<="000000000000001101000110";
t(1890)<="000000000000010001001000";
t(1891)<="000000000000010100111100";
t(1892)<="000000000000011000011100";
t(1893)<="000000000000011011100110";
t(1894)<="000000000000011110010101";
t(1895)<="000000000000100000101000";
t(1896)<="000000000000100010011100";
t(1897)<="000000000000100011101111";
t(1898)<="000000000000100100011110";
t(1899)<="000000000000100100101010";
t(1900)<="000000000000100100010001";
t(1901)<="000000000000100011010100";
t(1902)<="000000000000100001110011";
t(1903)<="000000000000011111110000";
t(1904)<="000000000000011101001011";
t(1905)<="000000000000011010001001";
t(1906)<="000000000000010110101001";
t(1907)<="000000000000010010110001";
t(1908)<="000000000000001110100011";
t(1909)<="000000000000001010000100";
t(1910)<="000000000000000101010110";
t(1911)<="000000000000000000100000";
t(1912)<="111111111111111111111111";
t(1913)<="111111111111111111111111";
t(1914)<="111111111111110001110011";
t(1915)<="111111111111101101000101";
t(1916)<="111111111111101000100101";
t(1917)<="111111111111100100011000";
t(1918)<="111111111111100000100001";
t(1919)<="111111111111011101000100";
t(1920)<="111111111111011010000101";
t(1921)<="111111111111010111100111";
t(1922)<="111111111111010101101101";
t(1923)<="111111111111010100011001";
t(1924)<="111111111111010011101100";
t(1925)<="111111111111010011101000";
t(1926)<="111111111111010100001110";
t(1927)<="111111111111010101011110";
t(1928)<="111111111111010111010110";
t(1929)<="111111111111011001110111";
t(1930)<="111111111111011100111101";
t(1931)<="111111111111100000101000";
t(1932)<="111111111111100100110100";
t(1933)<="111111111111101001011111";
t(1934)<="111111111111101110100011";
t(1935)<="111111111111111111111111";
t(1936)<="111111111111111111111111";
t(1937)<="111111111111111111111111";
t(1938)<="000000000000000101101011";
t(1939)<="000000000000001011110010";
t(1940)<="000000000000010001111000";
t(1941)<="000000000000010111110111";
t(1942)<="000000000000011101101010";
t(1943)<="000000000000100011001100";
t(1944)<="000000000000101000011000";
t(1945)<="000000000000101101001001";
t(1946)<="000000000000110001011011";
t(1947)<="000000000000110101001011";
t(1948)<="000000000000111000010011";
t(1949)<="000000000000111010110010";
t(1950)<="000000000000111100100011";
t(1951)<="000000000000111101100101";
t(1952)<="000000000000111101110111";
t(1953)<="000000000000111101010110";
t(1954)<="000000000000111100000010";
t(1955)<="000000000000111001111100";
t(1956)<="000000000000110111000011";
t(1957)<="000000000000110011011001";
t(1958)<="000000000000101110111111";
t(1959)<="000000000000101001110111";
t(1960)<="000000000000100100000100";
t(1961)<="000000000000011101101010";
t(1962)<="000000000000010110101010";
t(1963)<="000000000000001111001010";
t(1964)<="000000000000000111001110";
t(1965)<="111111111111111111111111";
t(1966)<="111111111111111111111111";
t(1967)<="111111111111101101011010";
t(1968)<="111111111111100100011011";
t(1969)<="111111111111011011010101";
t(1970)<="111111111111010010010011";
t(1971)<="111111111111001001010100";
t(1972)<="111111111111000000011101";
t(1973)<="111111111110110111111011";
t(1974)<="111111111110101111101001";
t(1975)<="111111111110100111101111";
t(1976)<="111111111110100000010001";
t(1977)<="111111111110011001010100";
t(1978)<="111111111110010010111000";
t(1979)<="111111111110001101000010";
t(1980)<="111111111110000111110010";
t(1981)<="111111111110000011001111";
t(1982)<="111111111101111111010111";
t(1983)<="111111111101111100001100";
t(1984)<="111111111101111001101100";
t(1985)<="111111111101110111111011";
t(1986)<="111111111101110110110110";
t(1987)<="111111111101110110100000";
t(1988)<="111111111101110110110100";
t(1989)<="111111111101110111110011";
t(1990)<="111111111101111001011001";
t(1991)<="111111111101111011100110";
t(1992)<="111111111101111110010110";
t(1993)<="111111111110000001101001";
t(1994)<="111111111110000101011001";
t(1995)<="111111111110001001100101";
t(1996)<="111111111110001110001001";
t(1997)<="111111111110010011000011";
t(1998)<="111111111110011000001101";
t(1999)<="111111111110011101100110";
t(2000)<="111111111110100011001001";
t(2001)<="111111111110101000110100";
t(2002)<="111111111110101110100100";
t(2003)<="111111111110110100010101";
t(2004)<="111111111110111010000101";
t(2005)<="111111111110111111110001";
t(2006)<="111111111111000101010110";
t(2007)<="111111111111001010110010";
t(2008)<="111111111111010000000010";
t(2009)<="111111111111010101000101";
t(2010)<="111111111111011001111001";
t(2011)<="111111111111011110011110";
t(2012)<="111111111111100010110000";
t(2013)<="111111111111100110110001";
t(2014)<="111111111111101010011100";
t(2015)<="111111111111101111000100";
t(2016)<="111111111111010010101011";
t(2017)<="111111111111111111111111";


        
    elsif (rising_edge(clk)) then
--------------------------------------------------------------------    
-----------------------------SENDING OUT ---------------------------    
--------------------------------------------------------------------       
        if(clk250k = '1') then   
		Load_On<='1';
        	a_s <= (others => '0');
        	b_s <= (others => '0');
        	c_s <= (others => '0');
        	d_s <= (others => '0');
        	e_s <= (others => '0');
		f_s <= (others => '0');
            	finished_sig <= '0';
           	finished<='0';
         	i<=0;
	elsif(finished_sig = '0' AND Load_On='0' AND GoOn='1') then
		if(i<N/6) then
			a_s <= a_s + (queue2multi(6*i)*t(6*i));
			b_s <= b_s + (queue2multi(6*i+1)*t(6*i+1));
			c_s <= c_s + (queue2multi(6*i+2)*t(6*i+2));
			d_s <= d_s + (queue2multi(6*i+3)*t(6*i+3));
			e_s <= e_s + (queue2multi(6*i+4)*t(6*i+4));
			f_s <= f_s + (queue2multi(6*i+5)*t(6*i+5));
			i <= i+1;
		else
			finished <= '1';
               		finished_sig <= '1';
                	y <= (a_s(2*width-2 downto width+11) + b_s(2*width-2 downto width+11) + c_s(2*width-2 downto width+11) + d_s(2*width-2 downto width+11) + e_s(2*width-2 downto width+11) + f_s(2*width-2 downto width+11));
                end if;
		
        end if;
--------------------------------------------------------------------    
-----------------------------READING IN ----------------------------    
--------------------------------------------------------------------  

	if (clk6M='1' ) then 
		pipe <= signed(x_sig)&pipe(0 to pipe'length-2);
	elsif(Load_On ='1') then
		for j in 0 to N-1 loop
             	   queue2multi(j)<= pipe(j);
         	end loop;
		GoOn<='1';  
		Load_On<='0';
	end if;

    end if;
end process;

end behaiv_arch;

