


-- This is a Linear phase FIR filter of type 1. Has N coeff. and N-1 inputs.
-- The filter is written generic so it is defined as;
--                            Width = number of bits
--                            N = number of tabs   
--			      M = Channel filter type, (to maximise the available space for multiplication)
-- Takes in, generic values width (nr. of bits), N number of tabs, x[n].
-- Sends out finihs signal, and y[n] (note double size, need to take the 12 last bits)
-- Authors: Jo³n Trausti
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Block_Filter_250 is
    generic(Width    :integer     :=12;
        N :integer    :=188);
    port(    reset:IN STD_LOGIC;
           clk:IN STD_LOGIC;
           clk250k:IN STD_LOGIC;
           clk4M:IN STD_LOGIC;
           x:IN signed(width-1-4 DOWNTO 0);
           y:OUT signed(WIDTH-1-4 DOWNTO 0);
           finished:OUT STD_LOGIC);
end Block_Filter_250;



architecture behaiv_arch of Block_Filter_250 is


-- New signals
signal i    :integer range 0 to N+3; --index for how many clkcykles the calculation have been running
signal finished_sig,GoOn,Load_On    :std_logic :='0';
signal y_s    :signed(2*width-1 downto 0);--temporary output
signal x_sig :signed(width-1 downto 0);

type a_pipe is array (0 to N-1) of signed(width-1 downto 0);
type a_queue2multi is array (0 to N-1) of signed(width-1 downto 0);
type a_tL is array (0 to N-1) of signed(width-1 downto 0);

signal pipe    		: a_pipe;
signal queue2multi	:a_queue2multi;
signal t		:a_tL;




-- Old signals



begin


x_sig(width-1 downto 4) <= x;
x_sig(3 downto 0) <= (others => '0');
process(clk,reset)
begin

    -- This will set all the x's to zero, resetting everything.
    -- so when the program start all values have zeros except for the coefficients
    if(reset='1') then
        i<=0;    -- reset the counter
        y_s <= (others => '0');
        y <= (others => '0');
        finished <= '0';
        finished_sig <= '1';
        for i in 0 to (N-1) loop
               pipe(i)<=(others=> '0');
               queue2multi(i)<=(others=> '0');
        end loop;
        

        -- here the coeff. comes in for ex.
t(0)<="0000000000001001";
        t(1)<="1111111111001001";
        t(2)<="1111111100010000";
        t(3)<="1111111001011010";
        t(4)<="1111111010011001";
        t(5)<="1111111111010010";
        t(6)<="0000000010111001";
        t(7)<="0000000001011100";
        t(8)<="1111111110010000";
        t(9)<="1111111110100010";
        t(10)<="0000000001001100";
        t(11)<="0000000001010110";
        t(12)<="1111111111000011";
        t(13)<="1111111110101111";
        t(14)<="0000000000110100";
        t(15)<="0000000001001011";
        t(16)<="1111111111001101";
        t(17)<="1111111110111000";
        t(18)<="0000000000110011";
        t(19)<="0000000001000101";
        t(20)<="1111111111001010";
        t(21)<="1111111110111011";
        t(22)<="0000000000111001";
        t(23)<="0000000001000011";
        t(24)<="1111111111000001";
        t(25)<="1111111110111100";
        t(26)<="0000000001000100";
        t(27)<="0000000001000011";
        t(28)<="1111111110110101";
        t(29)<="1111111110111100";
        t(30)<="0000000001010001";
        t(31)<="0000000001000011";
        t(32)<="1111111110100110";
        t(33)<="1111111110111100";
        t(34)<="0000000001100010";
        t(35)<="0000000001000011";
        t(36)<="1111111110010100";
        t(37)<="1111111110111101";
        t(38)<="0000000001110110";
        t(39)<="0000000001000000";
        t(40)<="1111111101111110";
        t(41)<="1111111111000000";
        t(42)<="0000000010001101";
        t(43)<="0000000000111100";
        t(44)<="1111111101100101";
        t(45)<="1111111111000110";
        t(46)<="0000000010101000";
        t(47)<="0000000000110101";
        t(48)<="1111111101001001";
        t(49)<="1111111111001111";
        t(50)<="0000000011000110";
        t(51)<="0000000000101010";
        t(52)<="1111111100100111";
        t(53)<="1111111111011101";
        t(54)<="0000000011101010";
        t(55)<="0000000000011001";
        t(56)<="1111111100000001";
        t(57)<="1111111111110000";
        t(58)<="0000000100010011";
        t(59)<="0000000000000010";
        t(60)<="1111111011010100";
        t(61)<="0000000000001100";
        t(62)<="0000000101000101";
        t(63)<="1111111111100001";
        t(64)<="1111111010011110";
        t(65)<="0000000000110011";
        t(66)<="0000000110000001";
        t(67)<="1111111110110010";
        t(68)<="1111111001011010";
        t(69)<="0000000001101011";
        t(70)<="0000000111001110";
        t(71)<="1111111101101111";
        t(72)<="1111111000000001";
        t(73)<="0000000010111110";
        t(74)<="0000001000111000";
        t(75)<="1111111100001000";
        t(76)<="1111110110000001";
        t(77)<="0000000101000001";
        t(78)<="0000001011011000";
        t(79)<="1111111001011011";
        t(80)<="1111110010101110";
        t(81)<="0000001000110000";
        t(82)<="0000001111111111";
        t(83)<="1111110011111011";
        t(84)<="1111101011101101";
        t(85)<="0000010001101111";
        t(86)<="0000011100010010";
        t(87)<="1111100010001100";
        t(88)<="1111001111000110";
        t(89)<="0001001001110011";
        t(90)<="0011101001011001";
        t(91)<="0011101001011001";
        t(92)<="0001001001110011";
        t(93)<="1111001111000110";
        t(94)<="1111100010001100";
        t(95)<="0000011100010010";
        t(96)<="0000010001101111";
        t(97)<="1111101011101101";
        t(98)<="1111110011111011";
        t(99)<="0000001111111111";
        t(100)<="0000001000110000";
        t(101)<="1111110010101110";
        t(102)<="1111111001011011";
        t(103)<="0000001011011000";
        t(104)<="0000000101000001";
        t(105)<="1111110110000001";
        t(106)<="1111111100001000";
        t(107)<="0000001000111000";
        t(108)<="0000000010111110";
        t(109)<="1111111000000001";
        t(110)<="1111111101101111";
        t(111)<="0000000111001110";
        t(112)<="0000000001101011";
        t(113)<="1111111001011010";
        t(114)<="1111111110110010";
        t(115)<="0000000110000001";
        t(116)<="0000000000110011";
        t(117)<="1111111010011110";
        t(118)<="1111111111100001";
        t(119)<="0000000101000101";
        t(120)<="0000000000001100";
        t(121)<="1111111011010100";
        t(122)<="0000000000000010";
        t(123)<="0000000100010011";
        t(124)<="1111111111110000";
        t(125)<="1111111100000001";
        t(126)<="0000000000011001";
        t(127)<="0000000011101010";
        t(128)<="1111111111011101";
        t(129)<="1111111100100111";
        t(130)<="0000000000101010";
        t(131)<="0000000011000110";
        t(132)<="1111111111001111";
        t(133)<="1111111101001001";
        t(134)<="0000000000110101";
        t(135)<="0000000010101000";
        t(136)<="1111111111000110";
        t(137)<="1111111101100101";
        t(138)<="0000000000111100";
        t(139)<="0000000010001101";
        t(140)<="1111111111000000";
        t(141)<="1111111101111110";
        t(142)<="0000000001000000";
        t(143)<="0000000001110110";
        t(144)<="1111111110111101";
        t(145)<="1111111110010100";
        t(146)<="0000000001000011";
        t(147)<="0000000001100010";
        t(148)<="1111111110111100";
        t(149)<="1111111110100110";
        t(150)<="0000000001000011";
        t(151)<="0000000001010001";
        t(152)<="1111111110111100";
        t(153)<="1111111110110101";
        t(154)<="0000000001000011";
        t(155)<="0000000001000100";
        t(156)<="1111111110111100";
        t(157)<="1111111111000001";
        t(158)<="0000000001000011";
        t(159)<="0000000000111001";
        t(160)<="1111111110111011";
        t(161)<="1111111111001010";
        t(162)<="0000000001000101";
        t(163)<="0000000000110011";
        t(164)<="1111111110111000";
        t(165)<="1111111111001101";
        t(166)<="0000000001001011";
        t(167)<="0000000000110100";
        t(168)<="1111111110101111";
        t(169)<="1111111111000011";
        t(170)<="0000000001010110";
        t(171)<="0000000001001100";
        t(172)<="1111111110100010";
        t(173)<="1111111110010000";
        t(174)<="0000000001011100";
        t(175)<="0000000010111001";
        t(176)<="1111111111010010";
        t(177)<="1111111010011001";
        t(178)<="1111111001011010";
        t(179)<="1111111100010000";
        t(180)<="1111111111001001";
        t(181)<="0000000000001001";




    elsif (rising_edge(clk)) then
--------------------------------------------------------------------    
-----------------------------SENDING OUT ---------------------------    
--------------------------------------------------------------------       
        if(clk250k = '1') then   
		Load_On<='1';
        	y_s <= (others => '0');
            	finished_sig <= '0';
           	finished<='0';
         	i<=0;
	elsif(finished_sig = '0' AND Load_On='0' AND GoOn='1') then
		if(i<N) then
			y_s <= y_s + (queue2multi(i)*t(i));
			i <= i+1;
		else
			finished <= '1';
                	finished_sig <= '1';
               		y <= y_s(2*width-2 downto width-1+4);
		end if;
		
        end if;
--------------------------------------------------------------------    
-----------------------------READING IN ----------------------------    
--------------------------------------------------------------------  

	if (clk4M='1' ) then 
		pipe <= signed(x_sig)&pipe(0 to pipe'length-2);
	elsif(Load_On ='1') then
		for j in 0 to N-1 loop
             	   queue2multi(j)<= pipe(j);
         	end loop;
		GoOn<='1';  
		Load_On<='0';
	end if;

    end if;
end process;

end behaiv_arch;
