


-- This is a Linear phase FIR filter of type 1. Has N coeff. and N-1 inputs.
-- The filter is written generic so it is defined as;
--                            Width = number of bits
--                            N = number of tabs   
--			      M = Channel filter type, (to maximise the available space for multiplication)
-- Takes in, generic values width (nr. of bits), N number of tabs, x[n].
-- Sends out finihs signal, and y[n] (note double size, need to take the 12 last bits)
-- Authors: Jo³n Trausti
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Block_Filter_250 is
    generic(Width    :integer     :=12;
        N :integer    :=188);
    port(    reset:IN STD_LOGIC;
           clk:IN STD_LOGIC;
           clk250k:IN STD_LOGIC;
           clk4M:IN STD_LOGIC;
           x:IN signed(width-1-4 DOWNTO 0);
           y:OUT signed(WIDTH-1-4 DOWNTO 0);
           finished:OUT STD_LOGIC);
end Block_Filter_250;



architecture behaiv_arch of Block_Filter_250 is


-- New signals
signal i    :integer range 0 to N+3; --index for how many clkcykles the calculation have been running
signal finished_sig,GoOn,Load_On    :std_logic :='0';
signal y_s    :signed(2*width-1 downto 0);--temporary output
signal x_sig :signed(width-1 downto 0);

type a_pipe is array (0 to N-1) of signed(width-1 downto 0);
type a_queue2multi is array (0 to N-1) of signed(width-1 downto 0);
type a_tL is array (0 to N-1) of signed(width-1 downto 0);

signal pipe    		: a_pipe;
signal queue2multi	:a_queue2multi;
signal t		:a_tL;




-- Old signals



begin


x_sig(width-1 downto 4) <= x;
x_sig(3 downto 0) <= (others => '0');
process(clk,reset)
begin

    -- This will set all the x's to zero, resetting everything.
    -- so when the program start all values have zeros except for the coefficients
    if(reset='1') then
        i<=0;    -- reset the counter
        y_s <= (others => '0');
        y <= (others => '0');
        finished <= '0';
        finished_sig <= '1';
        for i in 0 to (N-1) loop
               pipe(i)<=(others=> '0');
               queue2multi(i)<=(others=> '0');
        end loop;
        

        -- here the coeff. comes in for ex.
        t(0)<="1111111111101011";
        t(1)<="1111111101110110";
        t(2)<="1111111011000000";
        t(3)<="1111111001101010";
        t(4)<="1111111100001101";
        t(5)<="0000000000110111";
        t(6)<="0000000010111101";
        t(7)<="0000000000110001";
        t(8)<="1111111110000100";
        t(9)<="1111111110101111";
        t(10)<="0000000001001110";
        t(11)<="0000000001010111";
        t(12)<="1111111111001110";
        t(13)<="1111111110100111";
        t(14)<="0000000000011101";
        t(15)<="0000000001010111";
        t(16)<="1111111111110000";
        t(17)<="1111111110101001";
        t(18)<="0000000000000011";
        t(19)<="0000000001010110";
        t(20)<="0000000000000111";
        t(21)<="1111111110101001";
        t(22)<="1111111111101110";
        t(23)<="0000000001010111";
        t(24)<="0000000000011100";
        t(25)<="1111111110101000";
        t(26)<="1111111111011000";
        t(27)<="0000000001010110";
        t(28)<="0000000000110011";
        t(29)<="1111111110101010";
        t(30)<="1111111110111111";
        t(31)<="0000000001010011";
        t(32)<="0000000001001101";
        t(33)<="1111111110110000";
        t(34)<="1111111110100100";
        t(35)<="0000000001001001";
        t(36)<="0000000001101010";
        t(37)<="1111111110111101";
        t(38)<="1111111110000111";
        t(39)<="0000000000111000";
        t(40)<="0000000010000111";
        t(41)<="1111111111010010";
        t(42)<="1111111101101010";
        t(43)<="0000000000011111";
        t(44)<="0000000010100011";
        t(45)<="1111111111110000";
        t(46)<="1111111101001110";
        t(47)<="1111111111111011";
        t(48)<="0000000010111101";
        t(49)<="0000000000011001";
        t(50)<="1111111100110111";
        t(51)<="1111111111001101";
        t(52)<="0000000011010001";
        t(53)<="0000000001001110";
        t(54)<="1111111100100110";
        t(55)<="1111111110010011";
        t(56)<="0000000011011110";
        t(57)<="0000000010001110";
        t(58)<="1111111100011111";
        t(59)<="1111111101001100";
        t(60)<="0000000011011111";
        t(61)<="0000000011011100";
        t(62)<="1111111100100101";
        t(63)<="1111111011110111";
        t(64)<="0000000011010000";
        t(65)<="0000000100111001";
        t(66)<="1111111100111110";
        t(67)<="1111111010010000";
        t(68)<="0000000010101100";
        t(69)<="0000000110101001";
        t(70)<="1111111101110000";
        t(71)<="1111111000010101";
        t(72)<="0000000001101001";
        t(73)<="0000001000110100";
        t(74)<="1111111111001000";
        t(75)<="1111110101110101";
        t(76)<="1111111111110100";
        t(77)<="0000001011101111";
        t(78)<="0000000001100011";
        t(79)<="1111110010010011";
        t(80)<="1111111100100010";
        t(81)<="0000010000010001";
        t(82)<="0000000110001111";
        t(83)<="1111101100000010";
        t(84)<="1111110101010111";
        t(85)<="0000011001111110";
        t(86)<="0000010010110010";
        t(87)<="1111011001101000";
        t(88)<="1111011000011100";
        t(89)<="0001010010101010";
        t(90)<="0011100000010010";
        t(91)<="0011100000010010";
        t(92)<="0001010010101010";
        t(93)<="1111011000011100";
        t(94)<="1111011001101000";
        t(95)<="0000010010110010";
        t(96)<="0000011001111110";
        t(97)<="1111110101010111";
        t(98)<="1111101100000010";
        t(99)<="0000000110001111";
        t(100)<="0000010000010001";
        t(101)<="1111111100100010";
        t(102)<="1111110010010011";
        t(103)<="0000000001100011";
        t(104)<="0000001011101111";
        t(105)<="1111111111110100";
        t(106)<="1111110101110101";
        t(107)<="1111111111001000";
        t(108)<="0000001000110100";
        t(109)<="0000000001101001";
        t(110)<="1111111000010101";
        t(111)<="1111111101110000";
        t(112)<="0000000110101001";
        t(113)<="0000000010101100";
        t(114)<="1111111010010000";
        t(115)<="1111111100111110";
        t(116)<="0000000100111001";
        t(117)<="0000000011010000";
        t(118)<="1111111011110111";
        t(119)<="1111111100100101";
        t(120)<="0000000011011100";
        t(121)<="0000000011011111";
        t(122)<="1111111101001100";
        t(123)<="1111111100011111";
        t(124)<="0000000010001110";
        t(125)<="0000000011011110";
        t(126)<="1111111110010011";
        t(127)<="1111111100100110";
        t(128)<="0000000001001110";
        t(129)<="0000000011010001";
        t(130)<="1111111111001101";
        t(131)<="1111111100110111";
        t(132)<="0000000000011001";
        t(133)<="0000000010111101";
        t(134)<="1111111111111011";
        t(135)<="1111111101001110";
        t(136)<="1111111111110000";
        t(137)<="0000000010100011";
        t(138)<="0000000000011111";
        t(139)<="1111111101101010";
        t(140)<="1111111111010010";
        t(141)<="0000000010000111";
        t(142)<="0000000000111000";
        t(143)<="1111111110000111";
        t(144)<="1111111110111101";
        t(145)<="0000000001101010";
        t(146)<="0000000001001001";
        t(147)<="1111111110100100";
        t(148)<="1111111110110000";
        t(149)<="0000000001001101";
        t(150)<="0000000001010011";
        t(151)<="1111111110111111";
        t(152)<="1111111110101010";
        t(153)<="0000000000110011";
        t(154)<="0000000001010110";
        t(155)<="1111111111011000";
        t(156)<="1111111110101000";
        t(157)<="0000000000011100";
        t(158)<="0000000001010111";
        t(159)<="1111111111101110";
        t(160)<="1111111110101001";
        t(161)<="0000000000000111";
        t(162)<="0000000001010110";
        t(163)<="0000000000000011";
        t(164)<="1111111110101001";
        t(165)<="1111111111110000";
        t(166)<="0000000001010111";
        t(167)<="0000000000011101";
        t(168)<="1111111110100111";
        t(169)<="1111111111001110";
        t(170)<="0000000001010111";
        t(171)<="0000000001001110";
        t(172)<="1111111110101111";
        t(173)<="1111111110000100";
        t(174)<="0000000000110001";
        t(175)<="0000000010111101";
        t(176)<="0000000000110111";
        t(177)<="1111111100001101";
        t(178)<="1111111001101010";
        t(179)<="1111111011000000";
        t(180)<="1111111101110110";
        t(181)<="1111111111101011";



    elsif (rising_edge(clk)) then
--------------------------------------------------------------------    
-----------------------------SENDING OUT ---------------------------    
--------------------------------------------------------------------       
        if(clk250k = '1') then   
		Load_On<='1';
        	y_s <= (others => '0');
            	finished_sig <= '0';
           	finished<='0';
         	i<=0;
	elsif(finished_sig = '0' AND Load_On='0' AND GoOn='1') then
		if(i<N) then
			y_s <= y_s + (queue2multi(i)*t(i));
			i <= i+1;
		else
			finished <= '1';
                	finished_sig <= '1';
               		y <= y_s(2*width-2 downto width-1+4);
		end if;
		
        end if;
--------------------------------------------------------------------    
-----------------------------READING IN ----------------------------    
--------------------------------------------------------------------  

	if (clk4M='1' ) then 
		pipe <= signed(x_sig)&pipe(0 to pipe'length-2);
	elsif(Load_On ='1') then
		for j in 0 to N-1 loop
             	   queue2multi(j)<= pipe(j);
         	end loop;
		GoOn<='1';  
		Load_On<='0';
	end if;

    end if;
end process;

end behaiv_arch;
